module sort_pipe(
     input clk,
     input  [7:0] x_0, x_1, x_2, x_3, x_4, x_5, x_6, x_7, x_8, x_9, x_10, x_11, x_12, x_13, x_14, x_15, x_16, x_17, x_18, x_19, x_20, x_21, x_22, x_23, x_24, x_25, x_26, x_27, x_28, x_29, x_30, x_31, x_32, x_33, x_34, x_35, x_36, x_37, x_38, x_39, x_40, x_41, x_42, x_43, x_44, x_45, x_46, x_47, x_48, x_49, x_50, x_51, x_52, x_53, x_54, x_55, x_56, x_57, x_58, x_59, x_60, x_61, x_62, x_63, x_64, x_65, x_66, x_67, x_68, x_69, x_70, x_71, x_72, x_73, x_74, x_75, x_76, x_77, x_78, x_79, x_80, 
     output [7:0] median
);
reg[7:0] r0 [80:0];
reg[7:0] r1 [80:0];
reg[7:0] r2 [80:0];
reg[7:0] r3 [80:0];
reg[7:0] r4 [80:0];
reg[7:0] r5 [80:0];
reg[7:0] r6 [80:0];
reg[7:0] r7 [80:0];
reg[7:0] r8 [80:0];
reg[7:0] r9 [80:0];
reg[7:0] r10 [80:0];
reg[7:0] r11 [80:0];
reg[7:0] r12 [80:0];
reg[7:0] r13 [80:0];
reg[7:0] r14 [80:0];
reg[7:0] r15 [80:0];
reg[7:0] r16 [80:0];
reg[7:0] r17 [80:0];
reg[7:0] r18 [80:0];
reg[7:0] r19 [80:0];
reg[7:0] r20 [80:0];
reg[7:0] r21 [80:0];
reg[7:0] r22 [80:0];
reg[7:0] r23 [80:0];
reg[7:0] r24 [80:0];
reg[7:0] r25 [80:0];
reg[7:0] r26 [80:0];
reg[7:0] r27 [80:0];

//-------declaration layer:0----------
wire [7:0] cmp0_out0;
wire [7:0] cmp0_out1;
reg [7:0] cmp0_in0;
reg [7:0] cmp0_in1;

wire [7:0] cmp1_out0;
wire [7:0] cmp1_out1;
reg [7:0] cmp1_in0;
reg [7:0] cmp1_in1;

wire [7:0] cmp2_out0;
wire [7:0] cmp2_out1;
reg [7:0] cmp2_in0;
reg [7:0] cmp2_in1;

wire [7:0] cmp3_out0;
wire [7:0] cmp3_out1;
reg [7:0] cmp3_in0;
reg [7:0] cmp3_in1;

wire [7:0] cmp4_out0;
wire [7:0] cmp4_out1;
reg [7:0] cmp4_in0;
reg [7:0] cmp4_in1;

wire [7:0] cmp5_out0;
wire [7:0] cmp5_out1;
reg [7:0] cmp5_in0;
reg [7:0] cmp5_in1;

wire [7:0] cmp6_out0;
wire [7:0] cmp6_out1;
reg [7:0] cmp6_in0;
reg [7:0] cmp6_in1;

wire [7:0] cmp7_out0;
wire [7:0] cmp7_out1;
reg [7:0] cmp7_in0;
reg [7:0] cmp7_in1;

wire [7:0] cmp8_out0;
wire [7:0] cmp8_out1;
reg [7:0] cmp8_in0;
reg [7:0] cmp8_in1;

wire [7:0] cmp9_out0;
wire [7:0] cmp9_out1;
reg [7:0] cmp9_in0;
reg [7:0] cmp9_in1;

wire [7:0] cmp10_out0;
wire [7:0] cmp10_out1;
reg [7:0] cmp10_in0;
reg [7:0] cmp10_in1;

wire [7:0] cmp11_out0;
wire [7:0] cmp11_out1;
reg [7:0] cmp11_in0;
reg [7:0] cmp11_in1;

wire [7:0] cmp12_out0;
wire [7:0] cmp12_out1;
reg [7:0] cmp12_in0;
reg [7:0] cmp12_in1;

wire [7:0] cmp13_out0;
wire [7:0] cmp13_out1;
reg [7:0] cmp13_in0;
reg [7:0] cmp13_in1;

wire [7:0] cmp14_out0;
wire [7:0] cmp14_out1;
reg [7:0] cmp14_in0;
reg [7:0] cmp14_in1;

wire [7:0] cmp15_out0;
wire [7:0] cmp15_out1;
reg [7:0] cmp15_in0;
reg [7:0] cmp15_in1;

wire [7:0] cmp16_out0;
wire [7:0] cmp16_out1;
reg [7:0] cmp16_in0;
reg [7:0] cmp16_in1;

//-------declaration layer:1----------
wire [7:0] cmp17_out0;
wire [7:0] cmp17_out1;
reg [7:0] cmp17_in0;
reg [7:0] cmp17_in1;

wire [7:0] cmp18_out0;
wire [7:0] cmp18_out1;
reg [7:0] cmp18_in0;
reg [7:0] cmp18_in1;

wire [7:0] cmp19_out0;
wire [7:0] cmp19_out1;
reg [7:0] cmp19_in0;
reg [7:0] cmp19_in1;

wire [7:0] cmp20_out0;
wire [7:0] cmp20_out1;
reg [7:0] cmp20_in0;
reg [7:0] cmp20_in1;

wire [7:0] cmp21_out0;
wire [7:0] cmp21_out1;
reg [7:0] cmp21_in0;
reg [7:0] cmp21_in1;

wire [7:0] cmp22_out0;
wire [7:0] cmp22_out1;
reg [7:0] cmp22_in0;
reg [7:0] cmp22_in1;

wire [7:0] cmp23_out0;
wire [7:0] cmp23_out1;
reg [7:0] cmp23_in0;
reg [7:0] cmp23_in1;

wire [7:0] cmp24_out0;
wire [7:0] cmp24_out1;
reg [7:0] cmp24_in0;
reg [7:0] cmp24_in1;

wire [7:0] cmp25_out0;
wire [7:0] cmp25_out1;
reg [7:0] cmp25_in0;
reg [7:0] cmp25_in1;

wire [7:0] cmp26_out0;
wire [7:0] cmp26_out1;
reg [7:0] cmp26_in0;
reg [7:0] cmp26_in1;

wire [7:0] cmp27_out0;
wire [7:0] cmp27_out1;
reg [7:0] cmp27_in0;
reg [7:0] cmp27_in1;

wire [7:0] cmp28_out0;
wire [7:0] cmp28_out1;
reg [7:0] cmp28_in0;
reg [7:0] cmp28_in1;

wire [7:0] cmp29_out0;
wire [7:0] cmp29_out1;
reg [7:0] cmp29_in0;
reg [7:0] cmp29_in1;

wire [7:0] cmp30_out0;
wire [7:0] cmp30_out1;
reg [7:0] cmp30_in0;
reg [7:0] cmp30_in1;

wire [7:0] cmp31_out0;
wire [7:0] cmp31_out1;
reg [7:0] cmp31_in0;
reg [7:0] cmp31_in1;

wire [7:0] cmp32_out0;
wire [7:0] cmp32_out1;
reg [7:0] cmp32_in0;
reg [7:0] cmp32_in1;

wire [7:0] cmp33_out0;
wire [7:0] cmp33_out1;
reg [7:0] cmp33_in0;
reg [7:0] cmp33_in1;

wire [7:0] cmp34_out0;
wire [7:0] cmp34_out1;
reg [7:0] cmp34_in0;
reg [7:0] cmp34_in1;

wire [7:0] cmp35_out0;
wire [7:0] cmp35_out1;
reg [7:0] cmp35_in0;
reg [7:0] cmp35_in1;

wire [7:0] cmp36_out0;
wire [7:0] cmp36_out1;
reg [7:0] cmp36_in0;
reg [7:0] cmp36_in1;

wire [7:0] cmp37_out0;
wire [7:0] cmp37_out1;
reg [7:0] cmp37_in0;
reg [7:0] cmp37_in1;

wire [7:0] cmp38_out0;
wire [7:0] cmp38_out1;
reg [7:0] cmp38_in0;
reg [7:0] cmp38_in1;

wire [7:0] cmp39_out0;
wire [7:0] cmp39_out1;
reg [7:0] cmp39_in0;
reg [7:0] cmp39_in1;

wire [7:0] cmp40_out0;
wire [7:0] cmp40_out1;
reg [7:0] cmp40_in0;
reg [7:0] cmp40_in1;

wire [7:0] cmp41_out0;
wire [7:0] cmp41_out1;
reg [7:0] cmp41_in0;
reg [7:0] cmp41_in1;

wire [7:0] cmp42_out0;
wire [7:0] cmp42_out1;
reg [7:0] cmp42_in0;
reg [7:0] cmp42_in1;

wire [7:0] cmp43_out0;
wire [7:0] cmp43_out1;
reg [7:0] cmp43_in0;
reg [7:0] cmp43_in1;

wire [7:0] cmp44_out0;
wire [7:0] cmp44_out1;
reg [7:0] cmp44_in0;
reg [7:0] cmp44_in1;

wire [7:0] cmp45_out0;
wire [7:0] cmp45_out1;
reg [7:0] cmp45_in0;
reg [7:0] cmp45_in1;

wire [7:0] cmp46_out0;
wire [7:0] cmp46_out1;
reg [7:0] cmp46_in0;
reg [7:0] cmp46_in1;

wire [7:0] cmp47_out0;
wire [7:0] cmp47_out1;
reg [7:0] cmp47_in0;
reg [7:0] cmp47_in1;

wire [7:0] cmp48_out0;
wire [7:0] cmp48_out1;
reg [7:0] cmp48_in0;
reg [7:0] cmp48_in1;

//-------declaration layer:2----------
wire [7:0] cmp49_out0;
wire [7:0] cmp49_out1;
reg [7:0] cmp49_in0;
reg [7:0] cmp49_in1;

wire [7:0] cmp50_out0;
wire [7:0] cmp50_out1;
reg [7:0] cmp50_in0;
reg [7:0] cmp50_in1;

wire [7:0] cmp51_out0;
wire [7:0] cmp51_out1;
reg [7:0] cmp51_in0;
reg [7:0] cmp51_in1;

wire [7:0] cmp52_out0;
wire [7:0] cmp52_out1;
reg [7:0] cmp52_in0;
reg [7:0] cmp52_in1;

wire [7:0] cmp53_out0;
wire [7:0] cmp53_out1;
reg [7:0] cmp53_in0;
reg [7:0] cmp53_in1;

wire [7:0] cmp54_out0;
wire [7:0] cmp54_out1;
reg [7:0] cmp54_in0;
reg [7:0] cmp54_in1;

wire [7:0] cmp55_out0;
wire [7:0] cmp55_out1;
reg [7:0] cmp55_in0;
reg [7:0] cmp55_in1;

wire [7:0] cmp56_out0;
wire [7:0] cmp56_out1;
reg [7:0] cmp56_in0;
reg [7:0] cmp56_in1;

wire [7:0] cmp57_out0;
wire [7:0] cmp57_out1;
reg [7:0] cmp57_in0;
reg [7:0] cmp57_in1;

wire [7:0] cmp58_out0;
wire [7:0] cmp58_out1;
reg [7:0] cmp58_in0;
reg [7:0] cmp58_in1;

wire [7:0] cmp59_out0;
wire [7:0] cmp59_out1;
reg [7:0] cmp59_in0;
reg [7:0] cmp59_in1;

wire [7:0] cmp60_out0;
wire [7:0] cmp60_out1;
reg [7:0] cmp60_in0;
reg [7:0] cmp60_in1;

wire [7:0] cmp61_out0;
wire [7:0] cmp61_out1;
reg [7:0] cmp61_in0;
reg [7:0] cmp61_in1;

wire [7:0] cmp62_out0;
wire [7:0] cmp62_out1;
reg [7:0] cmp62_in0;
reg [7:0] cmp62_in1;

wire [7:0] cmp63_out0;
wire [7:0] cmp63_out1;
reg [7:0] cmp63_in0;
reg [7:0] cmp63_in1;

wire [7:0] cmp64_out0;
wire [7:0] cmp64_out1;
reg [7:0] cmp64_in0;
reg [7:0] cmp64_in1;

wire [7:0] cmp65_out0;
wire [7:0] cmp65_out1;
reg [7:0] cmp65_in0;
reg [7:0] cmp65_in1;

wire [7:0] cmp66_out0;
wire [7:0] cmp66_out1;
reg [7:0] cmp66_in0;
reg [7:0] cmp66_in1;

wire [7:0] cmp67_out0;
wire [7:0] cmp67_out1;
reg [7:0] cmp67_in0;
reg [7:0] cmp67_in1;

wire [7:0] cmp68_out0;
wire [7:0] cmp68_out1;
reg [7:0] cmp68_in0;
reg [7:0] cmp68_in1;

wire [7:0] cmp69_out0;
wire [7:0] cmp69_out1;
reg [7:0] cmp69_in0;
reg [7:0] cmp69_in1;

wire [7:0] cmp70_out0;
wire [7:0] cmp70_out1;
reg [7:0] cmp70_in0;
reg [7:0] cmp70_in1;

wire [7:0] cmp71_out0;
wire [7:0] cmp71_out1;
reg [7:0] cmp71_in0;
reg [7:0] cmp71_in1;

wire [7:0] cmp72_out0;
wire [7:0] cmp72_out1;
reg [7:0] cmp72_in0;
reg [7:0] cmp72_in1;

wire [7:0] cmp73_out0;
wire [7:0] cmp73_out1;
reg [7:0] cmp73_in0;
reg [7:0] cmp73_in1;

wire [7:0] cmp74_out0;
wire [7:0] cmp74_out1;
reg [7:0] cmp74_in0;
reg [7:0] cmp74_in1;

wire [7:0] cmp75_out0;
wire [7:0] cmp75_out1;
reg [7:0] cmp75_in0;
reg [7:0] cmp75_in1;

wire [7:0] cmp76_out0;
wire [7:0] cmp76_out1;
reg [7:0] cmp76_in0;
reg [7:0] cmp76_in1;

wire [7:0] cmp77_out0;
wire [7:0] cmp77_out1;
reg [7:0] cmp77_in0;
reg [7:0] cmp77_in1;

wire [7:0] cmp78_out0;
wire [7:0] cmp78_out1;
reg [7:0] cmp78_in0;
reg [7:0] cmp78_in1;

wire [7:0] cmp79_out0;
wire [7:0] cmp79_out1;
reg [7:0] cmp79_in0;
reg [7:0] cmp79_in1;

wire [7:0] cmp80_out0;
wire [7:0] cmp80_out1;
reg [7:0] cmp80_in0;
reg [7:0] cmp80_in1;

wire [7:0] cmp81_out0;
wire [7:0] cmp81_out1;
reg [7:0] cmp81_in0;
reg [7:0] cmp81_in1;

//-------declaration layer:3----------
wire [7:0] cmp82_out0;
wire [7:0] cmp82_out1;
reg [7:0] cmp82_in0;
reg [7:0] cmp82_in1;

wire [7:0] cmp83_out0;
wire [7:0] cmp83_out1;
reg [7:0] cmp83_in0;
reg [7:0] cmp83_in1;

wire [7:0] cmp84_out0;
wire [7:0] cmp84_out1;
reg [7:0] cmp84_in0;
reg [7:0] cmp84_in1;

wire [7:0] cmp85_out0;
wire [7:0] cmp85_out1;
reg [7:0] cmp85_in0;
reg [7:0] cmp85_in1;

wire [7:0] cmp86_out0;
wire [7:0] cmp86_out1;
reg [7:0] cmp86_in0;
reg [7:0] cmp86_in1;

wire [7:0] cmp87_out0;
wire [7:0] cmp87_out1;
reg [7:0] cmp87_in0;
reg [7:0] cmp87_in1;

wire [7:0] cmp88_out0;
wire [7:0] cmp88_out1;
reg [7:0] cmp88_in0;
reg [7:0] cmp88_in1;

wire [7:0] cmp89_out0;
wire [7:0] cmp89_out1;
reg [7:0] cmp89_in0;
reg [7:0] cmp89_in1;

wire [7:0] cmp90_out0;
wire [7:0] cmp90_out1;
reg [7:0] cmp90_in0;
reg [7:0] cmp90_in1;

wire [7:0] cmp91_out0;
wire [7:0] cmp91_out1;
reg [7:0] cmp91_in0;
reg [7:0] cmp91_in1;

wire [7:0] cmp92_out0;
wire [7:0] cmp92_out1;
reg [7:0] cmp92_in0;
reg [7:0] cmp92_in1;

wire [7:0] cmp93_out0;
wire [7:0] cmp93_out1;
reg [7:0] cmp93_in0;
reg [7:0] cmp93_in1;

wire [7:0] cmp94_out0;
wire [7:0] cmp94_out1;
reg [7:0] cmp94_in0;
reg [7:0] cmp94_in1;

wire [7:0] cmp95_out0;
wire [7:0] cmp95_out1;
reg [7:0] cmp95_in0;
reg [7:0] cmp95_in1;

wire [7:0] cmp96_out0;
wire [7:0] cmp96_out1;
reg [7:0] cmp96_in0;
reg [7:0] cmp96_in1;

wire [7:0] cmp97_out0;
wire [7:0] cmp97_out1;
reg [7:0] cmp97_in0;
reg [7:0] cmp97_in1;

wire [7:0] cmp98_out0;
wire [7:0] cmp98_out1;
reg [7:0] cmp98_in0;
reg [7:0] cmp98_in1;

//-------declaration layer:4----------
wire [7:0] cmp99_out0;
wire [7:0] cmp99_out1;
reg [7:0] cmp99_in0;
reg [7:0] cmp99_in1;

wire [7:0] cmp100_out0;
wire [7:0] cmp100_out1;
reg [7:0] cmp100_in0;
reg [7:0] cmp100_in1;

wire [7:0] cmp101_out0;
wire [7:0] cmp101_out1;
reg [7:0] cmp101_in0;
reg [7:0] cmp101_in1;

wire [7:0] cmp102_out0;
wire [7:0] cmp102_out1;
reg [7:0] cmp102_in0;
reg [7:0] cmp102_in1;

wire [7:0] cmp103_out0;
wire [7:0] cmp103_out1;
reg [7:0] cmp103_in0;
reg [7:0] cmp103_in1;

wire [7:0] cmp104_out0;
wire [7:0] cmp104_out1;
reg [7:0] cmp104_in0;
reg [7:0] cmp104_in1;

wire [7:0] cmp105_out0;
wire [7:0] cmp105_out1;
reg [7:0] cmp105_in0;
reg [7:0] cmp105_in1;

wire [7:0] cmp106_out0;
wire [7:0] cmp106_out1;
reg [7:0] cmp106_in0;
reg [7:0] cmp106_in1;

wire [7:0] cmp107_out0;
wire [7:0] cmp107_out1;
reg [7:0] cmp107_in0;
reg [7:0] cmp107_in1;

wire [7:0] cmp108_out0;
wire [7:0] cmp108_out1;
reg [7:0] cmp108_in0;
reg [7:0] cmp108_in1;

wire [7:0] cmp109_out0;
wire [7:0] cmp109_out1;
reg [7:0] cmp109_in0;
reg [7:0] cmp109_in1;

wire [7:0] cmp110_out0;
wire [7:0] cmp110_out1;
reg [7:0] cmp110_in0;
reg [7:0] cmp110_in1;

wire [7:0] cmp111_out0;
wire [7:0] cmp111_out1;
reg [7:0] cmp111_in0;
reg [7:0] cmp111_in1;

wire [7:0] cmp112_out0;
wire [7:0] cmp112_out1;
reg [7:0] cmp112_in0;
reg [7:0] cmp112_in1;

wire [7:0] cmp113_out0;
wire [7:0] cmp113_out1;
reg [7:0] cmp113_in0;
reg [7:0] cmp113_in1;

wire [7:0] cmp114_out0;
wire [7:0] cmp114_out1;
reg [7:0] cmp114_in0;
reg [7:0] cmp114_in1;

//-------declaration layer:5----------
wire [7:0] cmp115_out0;
wire [7:0] cmp115_out1;
reg [7:0] cmp115_in0;
reg [7:0] cmp115_in1;

wire [7:0] cmp116_out0;
wire [7:0] cmp116_out1;
reg [7:0] cmp116_in0;
reg [7:0] cmp116_in1;

wire [7:0] cmp117_out0;
wire [7:0] cmp117_out1;
reg [7:0] cmp117_in0;
reg [7:0] cmp117_in1;

wire [7:0] cmp118_out0;
wire [7:0] cmp118_out1;
reg [7:0] cmp118_in0;
reg [7:0] cmp118_in1;

wire [7:0] cmp119_out0;
wire [7:0] cmp119_out1;
reg [7:0] cmp119_in0;
reg [7:0] cmp119_in1;

wire [7:0] cmp120_out0;
wire [7:0] cmp120_out1;
reg [7:0] cmp120_in0;
reg [7:0] cmp120_in1;

wire [7:0] cmp121_out0;
wire [7:0] cmp121_out1;
reg [7:0] cmp121_in0;
reg [7:0] cmp121_in1;

wire [7:0] cmp122_out0;
wire [7:0] cmp122_out1;
reg [7:0] cmp122_in0;
reg [7:0] cmp122_in1;

wire [7:0] cmp123_out0;
wire [7:0] cmp123_out1;
reg [7:0] cmp123_in0;
reg [7:0] cmp123_in1;

wire [7:0] cmp124_out0;
wire [7:0] cmp124_out1;
reg [7:0] cmp124_in0;
reg [7:0] cmp124_in1;

wire [7:0] cmp125_out0;
wire [7:0] cmp125_out1;
reg [7:0] cmp125_in0;
reg [7:0] cmp125_in1;

wire [7:0] cmp126_out0;
wire [7:0] cmp126_out1;
reg [7:0] cmp126_in0;
reg [7:0] cmp126_in1;

wire [7:0] cmp127_out0;
wire [7:0] cmp127_out1;
reg [7:0] cmp127_in0;
reg [7:0] cmp127_in1;

wire [7:0] cmp128_out0;
wire [7:0] cmp128_out1;
reg [7:0] cmp128_in0;
reg [7:0] cmp128_in1;

wire [7:0] cmp129_out0;
wire [7:0] cmp129_out1;
reg [7:0] cmp129_in0;
reg [7:0] cmp129_in1;

wire [7:0] cmp130_out0;
wire [7:0] cmp130_out1;
reg [7:0] cmp130_in0;
reg [7:0] cmp130_in1;

wire [7:0] cmp131_out0;
wire [7:0] cmp131_out1;
reg [7:0] cmp131_in0;
reg [7:0] cmp131_in1;

wire [7:0] cmp132_out0;
wire [7:0] cmp132_out1;
reg [7:0] cmp132_in0;
reg [7:0] cmp132_in1;

wire [7:0] cmp133_out0;
wire [7:0] cmp133_out1;
reg [7:0] cmp133_in0;
reg [7:0] cmp133_in1;

wire [7:0] cmp134_out0;
wire [7:0] cmp134_out1;
reg [7:0] cmp134_in0;
reg [7:0] cmp134_in1;

wire [7:0] cmp135_out0;
wire [7:0] cmp135_out1;
reg [7:0] cmp135_in0;
reg [7:0] cmp135_in1;

wire [7:0] cmp136_out0;
wire [7:0] cmp136_out1;
reg [7:0] cmp136_in0;
reg [7:0] cmp136_in1;

wire [7:0] cmp137_out0;
wire [7:0] cmp137_out1;
reg [7:0] cmp137_in0;
reg [7:0] cmp137_in1;

wire [7:0] cmp138_out0;
wire [7:0] cmp138_out1;
reg [7:0] cmp138_in0;
reg [7:0] cmp138_in1;

wire [7:0] cmp139_out0;
wire [7:0] cmp139_out1;
reg [7:0] cmp139_in0;
reg [7:0] cmp139_in1;

wire [7:0] cmp140_out0;
wire [7:0] cmp140_out1;
reg [7:0] cmp140_in0;
reg [7:0] cmp140_in1;

wire [7:0] cmp141_out0;
wire [7:0] cmp141_out1;
reg [7:0] cmp141_in0;
reg [7:0] cmp141_in1;

wire [7:0] cmp142_out0;
wire [7:0] cmp142_out1;
reg [7:0] cmp142_in0;
reg [7:0] cmp142_in1;

wire [7:0] cmp143_out0;
wire [7:0] cmp143_out1;
reg [7:0] cmp143_in0;
reg [7:0] cmp143_in1;

wire [7:0] cmp144_out0;
wire [7:0] cmp144_out1;
reg [7:0] cmp144_in0;
reg [7:0] cmp144_in1;

wire [7:0] cmp145_out0;
wire [7:0] cmp145_out1;
reg [7:0] cmp145_in0;
reg [7:0] cmp145_in1;

wire [7:0] cmp146_out0;
wire [7:0] cmp146_out1;
reg [7:0] cmp146_in0;
reg [7:0] cmp146_in1;

wire [7:0] cmp147_out0;
wire [7:0] cmp147_out1;
reg [7:0] cmp147_in0;
reg [7:0] cmp147_in1;

wire [7:0] cmp148_out0;
wire [7:0] cmp148_out1;
reg [7:0] cmp148_in0;
reg [7:0] cmp148_in1;

wire [7:0] cmp149_out0;
wire [7:0] cmp149_out1;
reg [7:0] cmp149_in0;
reg [7:0] cmp149_in1;

wire [7:0] cmp150_out0;
wire [7:0] cmp150_out1;
reg [7:0] cmp150_in0;
reg [7:0] cmp150_in1;

wire [7:0] cmp151_out0;
wire [7:0] cmp151_out1;
reg [7:0] cmp151_in0;
reg [7:0] cmp151_in1;

wire [7:0] cmp152_out0;
wire [7:0] cmp152_out1;
reg [7:0] cmp152_in0;
reg [7:0] cmp152_in1;

wire [7:0] cmp153_out0;
wire [7:0] cmp153_out1;
reg [7:0] cmp153_in0;
reg [7:0] cmp153_in1;

wire [7:0] cmp154_out0;
wire [7:0] cmp154_out1;
reg [7:0] cmp154_in0;
reg [7:0] cmp154_in1;

//-------declaration layer:6----------
wire [7:0] cmp155_out0;
wire [7:0] cmp155_out1;
reg [7:0] cmp155_in0;
reg [7:0] cmp155_in1;

wire [7:0] cmp156_out0;
wire [7:0] cmp156_out1;
reg [7:0] cmp156_in0;
reg [7:0] cmp156_in1;

wire [7:0] cmp157_out0;
wire [7:0] cmp157_out1;
reg [7:0] cmp157_in0;
reg [7:0] cmp157_in1;

wire [7:0] cmp158_out0;
wire [7:0] cmp158_out1;
reg [7:0] cmp158_in0;
reg [7:0] cmp158_in1;

wire [7:0] cmp159_out0;
wire [7:0] cmp159_out1;
reg [7:0] cmp159_in0;
reg [7:0] cmp159_in1;

wire [7:0] cmp160_out0;
wire [7:0] cmp160_out1;
reg [7:0] cmp160_in0;
reg [7:0] cmp160_in1;

wire [7:0] cmp161_out0;
wire [7:0] cmp161_out1;
reg [7:0] cmp161_in0;
reg [7:0] cmp161_in1;

wire [7:0] cmp162_out0;
wire [7:0] cmp162_out1;
reg [7:0] cmp162_in0;
reg [7:0] cmp162_in1;

wire [7:0] cmp163_out0;
wire [7:0] cmp163_out1;
reg [7:0] cmp163_in0;
reg [7:0] cmp163_in1;

wire [7:0] cmp164_out0;
wire [7:0] cmp164_out1;
reg [7:0] cmp164_in0;
reg [7:0] cmp164_in1;

wire [7:0] cmp165_out0;
wire [7:0] cmp165_out1;
reg [7:0] cmp165_in0;
reg [7:0] cmp165_in1;

wire [7:0] cmp166_out0;
wire [7:0] cmp166_out1;
reg [7:0] cmp166_in0;
reg [7:0] cmp166_in1;

wire [7:0] cmp167_out0;
wire [7:0] cmp167_out1;
reg [7:0] cmp167_in0;
reg [7:0] cmp167_in1;

wire [7:0] cmp168_out0;
wire [7:0] cmp168_out1;
reg [7:0] cmp168_in0;
reg [7:0] cmp168_in1;

wire [7:0] cmp169_out0;
wire [7:0] cmp169_out1;
reg [7:0] cmp169_in0;
reg [7:0] cmp169_in1;

wire [7:0] cmp170_out0;
wire [7:0] cmp170_out1;
reg [7:0] cmp170_in0;
reg [7:0] cmp170_in1;

wire [7:0] cmp171_out0;
wire [7:0] cmp171_out1;
reg [7:0] cmp171_in0;
reg [7:0] cmp171_in1;

wire [7:0] cmp172_out0;
wire [7:0] cmp172_out1;
reg [7:0] cmp172_in0;
reg [7:0] cmp172_in1;

wire [7:0] cmp173_out0;
wire [7:0] cmp173_out1;
reg [7:0] cmp173_in0;
reg [7:0] cmp173_in1;

wire [7:0] cmp174_out0;
wire [7:0] cmp174_out1;
reg [7:0] cmp174_in0;
reg [7:0] cmp174_in1;

wire [7:0] cmp175_out0;
wire [7:0] cmp175_out1;
reg [7:0] cmp175_in0;
reg [7:0] cmp175_in1;

wire [7:0] cmp176_out0;
wire [7:0] cmp176_out1;
reg [7:0] cmp176_in0;
reg [7:0] cmp176_in1;

wire [7:0] cmp177_out0;
wire [7:0] cmp177_out1;
reg [7:0] cmp177_in0;
reg [7:0] cmp177_in1;

wire [7:0] cmp178_out0;
wire [7:0] cmp178_out1;
reg [7:0] cmp178_in0;
reg [7:0] cmp178_in1;

wire [7:0] cmp179_out0;
wire [7:0] cmp179_out1;
reg [7:0] cmp179_in0;
reg [7:0] cmp179_in1;

wire [7:0] cmp180_out0;
wire [7:0] cmp180_out1;
reg [7:0] cmp180_in0;
reg [7:0] cmp180_in1;

wire [7:0] cmp181_out0;
wire [7:0] cmp181_out1;
reg [7:0] cmp181_in0;
reg [7:0] cmp181_in1;

wire [7:0] cmp182_out0;
wire [7:0] cmp182_out1;
reg [7:0] cmp182_in0;
reg [7:0] cmp182_in1;

wire [7:0] cmp183_out0;
wire [7:0] cmp183_out1;
reg [7:0] cmp183_in0;
reg [7:0] cmp183_in1;

wire [7:0] cmp184_out0;
wire [7:0] cmp184_out1;
reg [7:0] cmp184_in0;
reg [7:0] cmp184_in1;

wire [7:0] cmp185_out0;
wire [7:0] cmp185_out1;
reg [7:0] cmp185_in0;
reg [7:0] cmp185_in1;

wire [7:0] cmp186_out0;
wire [7:0] cmp186_out1;
reg [7:0] cmp186_in0;
reg [7:0] cmp186_in1;

//-------declaration layer:7----------
wire [7:0] cmp187_out0;
wire [7:0] cmp187_out1;
reg [7:0] cmp187_in0;
reg [7:0] cmp187_in1;

wire [7:0] cmp188_out0;
wire [7:0] cmp188_out1;
reg [7:0] cmp188_in0;
reg [7:0] cmp188_in1;

wire [7:0] cmp189_out0;
wire [7:0] cmp189_out1;
reg [7:0] cmp189_in0;
reg [7:0] cmp189_in1;

wire [7:0] cmp190_out0;
wire [7:0] cmp190_out1;
reg [7:0] cmp190_in0;
reg [7:0] cmp190_in1;

wire [7:0] cmp191_out0;
wire [7:0] cmp191_out1;
reg [7:0] cmp191_in0;
reg [7:0] cmp191_in1;

wire [7:0] cmp192_out0;
wire [7:0] cmp192_out1;
reg [7:0] cmp192_in0;
reg [7:0] cmp192_in1;

wire [7:0] cmp193_out0;
wire [7:0] cmp193_out1;
reg [7:0] cmp193_in0;
reg [7:0] cmp193_in1;

wire [7:0] cmp194_out0;
wire [7:0] cmp194_out1;
reg [7:0] cmp194_in0;
reg [7:0] cmp194_in1;

wire [7:0] cmp195_out0;
wire [7:0] cmp195_out1;
reg [7:0] cmp195_in0;
reg [7:0] cmp195_in1;

//-------declaration layer:8----------
wire [7:0] cmp196_out0;
wire [7:0] cmp196_out1;
reg [7:0] cmp196_in0;
reg [7:0] cmp196_in1;

wire [7:0] cmp197_out0;
wire [7:0] cmp197_out1;
reg [7:0] cmp197_in0;
reg [7:0] cmp197_in1;

wire [7:0] cmp198_out0;
wire [7:0] cmp198_out1;
reg [7:0] cmp198_in0;
reg [7:0] cmp198_in1;

wire [7:0] cmp199_out0;
wire [7:0] cmp199_out1;
reg [7:0] cmp199_in0;
reg [7:0] cmp199_in1;

wire [7:0] cmp200_out0;
wire [7:0] cmp200_out1;
reg [7:0] cmp200_in0;
reg [7:0] cmp200_in1;

wire [7:0] cmp201_out0;
wire [7:0] cmp201_out1;
reg [7:0] cmp201_in0;
reg [7:0] cmp201_in1;

wire [7:0] cmp202_out0;
wire [7:0] cmp202_out1;
reg [7:0] cmp202_in0;
reg [7:0] cmp202_in1;

wire [7:0] cmp203_out0;
wire [7:0] cmp203_out1;
reg [7:0] cmp203_in0;
reg [7:0] cmp203_in1;

wire [7:0] cmp204_out0;
wire [7:0] cmp204_out1;
reg [7:0] cmp204_in0;
reg [7:0] cmp204_in1;

wire [7:0] cmp205_out0;
wire [7:0] cmp205_out1;
reg [7:0] cmp205_in0;
reg [7:0] cmp205_in1;

wire [7:0] cmp206_out0;
wire [7:0] cmp206_out1;
reg [7:0] cmp206_in0;
reg [7:0] cmp206_in1;

wire [7:0] cmp207_out0;
wire [7:0] cmp207_out1;
reg [7:0] cmp207_in0;
reg [7:0] cmp207_in1;

wire [7:0] cmp208_out0;
wire [7:0] cmp208_out1;
reg [7:0] cmp208_in0;
reg [7:0] cmp208_in1;

wire [7:0] cmp209_out0;
wire [7:0] cmp209_out1;
reg [7:0] cmp209_in0;
reg [7:0] cmp209_in1;

wire [7:0] cmp210_out0;
wire [7:0] cmp210_out1;
reg [7:0] cmp210_in0;
reg [7:0] cmp210_in1;

wire [7:0] cmp211_out0;
wire [7:0] cmp211_out1;
reg [7:0] cmp211_in0;
reg [7:0] cmp211_in1;

wire [7:0] cmp212_out0;
wire [7:0] cmp212_out1;
reg [7:0] cmp212_in0;
reg [7:0] cmp212_in1;

wire [7:0] cmp213_out0;
wire [7:0] cmp213_out1;
reg [7:0] cmp213_in0;
reg [7:0] cmp213_in1;

wire [7:0] cmp214_out0;
wire [7:0] cmp214_out1;
reg [7:0] cmp214_in0;
reg [7:0] cmp214_in1;

wire [7:0] cmp215_out0;
wire [7:0] cmp215_out1;
reg [7:0] cmp215_in0;
reg [7:0] cmp215_in1;

wire [7:0] cmp216_out0;
wire [7:0] cmp216_out1;
reg [7:0] cmp216_in0;
reg [7:0] cmp216_in1;

wire [7:0] cmp217_out0;
wire [7:0] cmp217_out1;
reg [7:0] cmp217_in0;
reg [7:0] cmp217_in1;

wire [7:0] cmp218_out0;
wire [7:0] cmp218_out1;
reg [7:0] cmp218_in0;
reg [7:0] cmp218_in1;

wire [7:0] cmp219_out0;
wire [7:0] cmp219_out1;
reg [7:0] cmp219_in0;
reg [7:0] cmp219_in1;

wire [7:0] cmp220_out0;
wire [7:0] cmp220_out1;
reg [7:0] cmp220_in0;
reg [7:0] cmp220_in1;

//-------declaration layer:9----------
wire [7:0] cmp221_out0;
wire [7:0] cmp221_out1;
reg [7:0] cmp221_in0;
reg [7:0] cmp221_in1;

wire [7:0] cmp222_out0;
wire [7:0] cmp222_out1;
reg [7:0] cmp222_in0;
reg [7:0] cmp222_in1;

wire [7:0] cmp223_out0;
wire [7:0] cmp223_out1;
reg [7:0] cmp223_in0;
reg [7:0] cmp223_in1;

wire [7:0] cmp224_out0;
wire [7:0] cmp224_out1;
reg [7:0] cmp224_in0;
reg [7:0] cmp224_in1;

wire [7:0] cmp225_out0;
wire [7:0] cmp225_out1;
reg [7:0] cmp225_in0;
reg [7:0] cmp225_in1;

wire [7:0] cmp226_out0;
wire [7:0] cmp226_out1;
reg [7:0] cmp226_in0;
reg [7:0] cmp226_in1;

wire [7:0] cmp227_out0;
wire [7:0] cmp227_out1;
reg [7:0] cmp227_in0;
reg [7:0] cmp227_in1;

wire [7:0] cmp228_out0;
wire [7:0] cmp228_out1;
reg [7:0] cmp228_in0;
reg [7:0] cmp228_in1;

wire [7:0] cmp229_out0;
wire [7:0] cmp229_out1;
reg [7:0] cmp229_in0;
reg [7:0] cmp229_in1;

wire [7:0] cmp230_out0;
wire [7:0] cmp230_out1;
reg [7:0] cmp230_in0;
reg [7:0] cmp230_in1;

wire [7:0] cmp231_out0;
wire [7:0] cmp231_out1;
reg [7:0] cmp231_in0;
reg [7:0] cmp231_in1;

wire [7:0] cmp232_out0;
wire [7:0] cmp232_out1;
reg [7:0] cmp232_in0;
reg [7:0] cmp232_in1;

wire [7:0] cmp233_out0;
wire [7:0] cmp233_out1;
reg [7:0] cmp233_in0;
reg [7:0] cmp233_in1;

wire [7:0] cmp234_out0;
wire [7:0] cmp234_out1;
reg [7:0] cmp234_in0;
reg [7:0] cmp234_in1;

wire [7:0] cmp235_out0;
wire [7:0] cmp235_out1;
reg [7:0] cmp235_in0;
reg [7:0] cmp235_in1;

wire [7:0] cmp236_out0;
wire [7:0] cmp236_out1;
reg [7:0] cmp236_in0;
reg [7:0] cmp236_in1;

wire [7:0] cmp237_out0;
wire [7:0] cmp237_out1;
reg [7:0] cmp237_in0;
reg [7:0] cmp237_in1;

wire [7:0] cmp238_out0;
wire [7:0] cmp238_out1;
reg [7:0] cmp238_in0;
reg [7:0] cmp238_in1;

wire [7:0] cmp239_out0;
wire [7:0] cmp239_out1;
reg [7:0] cmp239_in0;
reg [7:0] cmp239_in1;

wire [7:0] cmp240_out0;
wire [7:0] cmp240_out1;
reg [7:0] cmp240_in0;
reg [7:0] cmp240_in1;

wire [7:0] cmp241_out0;
wire [7:0] cmp241_out1;
reg [7:0] cmp241_in0;
reg [7:0] cmp241_in1;

wire [7:0] cmp242_out0;
wire [7:0] cmp242_out1;
reg [7:0] cmp242_in0;
reg [7:0] cmp242_in1;

wire [7:0] cmp243_out0;
wire [7:0] cmp243_out1;
reg [7:0] cmp243_in0;
reg [7:0] cmp243_in1;

wire [7:0] cmp244_out0;
wire [7:0] cmp244_out1;
reg [7:0] cmp244_in0;
reg [7:0] cmp244_in1;

wire [7:0] cmp245_out0;
wire [7:0] cmp245_out1;
reg [7:0] cmp245_in0;
reg [7:0] cmp245_in1;

wire [7:0] cmp246_out0;
wire [7:0] cmp246_out1;
reg [7:0] cmp246_in0;
reg [7:0] cmp246_in1;

wire [7:0] cmp247_out0;
wire [7:0] cmp247_out1;
reg [7:0] cmp247_in0;
reg [7:0] cmp247_in1;

wire [7:0] cmp248_out0;
wire [7:0] cmp248_out1;
reg [7:0] cmp248_in0;
reg [7:0] cmp248_in1;

wire [7:0] cmp249_out0;
wire [7:0] cmp249_out1;
reg [7:0] cmp249_in0;
reg [7:0] cmp249_in1;

wire [7:0] cmp250_out0;
wire [7:0] cmp250_out1;
reg [7:0] cmp250_in0;
reg [7:0] cmp250_in1;

wire [7:0] cmp251_out0;
wire [7:0] cmp251_out1;
reg [7:0] cmp251_in0;
reg [7:0] cmp251_in1;

wire [7:0] cmp252_out0;
wire [7:0] cmp252_out1;
reg [7:0] cmp252_in0;
reg [7:0] cmp252_in1;

wire [7:0] cmp253_out0;
wire [7:0] cmp253_out1;
reg [7:0] cmp253_in0;
reg [7:0] cmp253_in1;

wire [7:0] cmp254_out0;
wire [7:0] cmp254_out1;
reg [7:0] cmp254_in0;
reg [7:0] cmp254_in1;

wire [7:0] cmp255_out0;
wire [7:0] cmp255_out1;
reg [7:0] cmp255_in0;
reg [7:0] cmp255_in1;

wire [7:0] cmp256_out0;
wire [7:0] cmp256_out1;
reg [7:0] cmp256_in0;
reg [7:0] cmp256_in1;

wire [7:0] cmp257_out0;
wire [7:0] cmp257_out1;
reg [7:0] cmp257_in0;
reg [7:0] cmp257_in1;

//-------declaration layer:10----------
wire [7:0] cmp258_out0;
wire [7:0] cmp258_out1;
reg [7:0] cmp258_in0;
reg [7:0] cmp258_in1;

wire [7:0] cmp259_out0;
wire [7:0] cmp259_out1;
reg [7:0] cmp259_in0;
reg [7:0] cmp259_in1;

wire [7:0] cmp260_out0;
wire [7:0] cmp260_out1;
reg [7:0] cmp260_in0;
reg [7:0] cmp260_in1;

wire [7:0] cmp261_out0;
wire [7:0] cmp261_out1;
reg [7:0] cmp261_in0;
reg [7:0] cmp261_in1;

wire [7:0] cmp262_out0;
wire [7:0] cmp262_out1;
reg [7:0] cmp262_in0;
reg [7:0] cmp262_in1;

wire [7:0] cmp263_out0;
wire [7:0] cmp263_out1;
reg [7:0] cmp263_in0;
reg [7:0] cmp263_in1;

wire [7:0] cmp264_out0;
wire [7:0] cmp264_out1;
reg [7:0] cmp264_in0;
reg [7:0] cmp264_in1;

wire [7:0] cmp265_out0;
wire [7:0] cmp265_out1;
reg [7:0] cmp265_in0;
reg [7:0] cmp265_in1;

wire [7:0] cmp266_out0;
wire [7:0] cmp266_out1;
reg [7:0] cmp266_in0;
reg [7:0] cmp266_in1;

wire [7:0] cmp267_out0;
wire [7:0] cmp267_out1;
reg [7:0] cmp267_in0;
reg [7:0] cmp267_in1;

wire [7:0] cmp268_out0;
wire [7:0] cmp268_out1;
reg [7:0] cmp268_in0;
reg [7:0] cmp268_in1;

wire [7:0] cmp269_out0;
wire [7:0] cmp269_out1;
reg [7:0] cmp269_in0;
reg [7:0] cmp269_in1;

wire [7:0] cmp270_out0;
wire [7:0] cmp270_out1;
reg [7:0] cmp270_in0;
reg [7:0] cmp270_in1;

wire [7:0] cmp271_out0;
wire [7:0] cmp271_out1;
reg [7:0] cmp271_in0;
reg [7:0] cmp271_in1;

wire [7:0] cmp272_out0;
wire [7:0] cmp272_out1;
reg [7:0] cmp272_in0;
reg [7:0] cmp272_in1;

wire [7:0] cmp273_out0;
wire [7:0] cmp273_out1;
reg [7:0] cmp273_in0;
reg [7:0] cmp273_in1;

wire [7:0] cmp274_out0;
wire [7:0] cmp274_out1;
reg [7:0] cmp274_in0;
reg [7:0] cmp274_in1;

wire [7:0] cmp275_out0;
wire [7:0] cmp275_out1;
reg [7:0] cmp275_in0;
reg [7:0] cmp275_in1;

wire [7:0] cmp276_out0;
wire [7:0] cmp276_out1;
reg [7:0] cmp276_in0;
reg [7:0] cmp276_in1;

wire [7:0] cmp277_out0;
wire [7:0] cmp277_out1;
reg [7:0] cmp277_in0;
reg [7:0] cmp277_in1;

wire [7:0] cmp278_out0;
wire [7:0] cmp278_out1;
reg [7:0] cmp278_in0;
reg [7:0] cmp278_in1;

wire [7:0] cmp279_out0;
wire [7:0] cmp279_out1;
reg [7:0] cmp279_in0;
reg [7:0] cmp279_in1;

wire [7:0] cmp280_out0;
wire [7:0] cmp280_out1;
reg [7:0] cmp280_in0;
reg [7:0] cmp280_in1;

wire [7:0] cmp281_out0;
wire [7:0] cmp281_out1;
reg [7:0] cmp281_in0;
reg [7:0] cmp281_in1;

wire [7:0] cmp282_out0;
wire [7:0] cmp282_out1;
reg [7:0] cmp282_in0;
reg [7:0] cmp282_in1;

wire [7:0] cmp283_out0;
wire [7:0] cmp283_out1;
reg [7:0] cmp283_in0;
reg [7:0] cmp283_in1;

wire [7:0] cmp284_out0;
wire [7:0] cmp284_out1;
reg [7:0] cmp284_in0;
reg [7:0] cmp284_in1;

wire [7:0] cmp285_out0;
wire [7:0] cmp285_out1;
reg [7:0] cmp285_in0;
reg [7:0] cmp285_in1;

wire [7:0] cmp286_out0;
wire [7:0] cmp286_out1;
reg [7:0] cmp286_in0;
reg [7:0] cmp286_in1;

wire [7:0] cmp287_out0;
wire [7:0] cmp287_out1;
reg [7:0] cmp287_in0;
reg [7:0] cmp287_in1;

wire [7:0] cmp288_out0;
wire [7:0] cmp288_out1;
reg [7:0] cmp288_in0;
reg [7:0] cmp288_in1;

wire [7:0] cmp289_out0;
wire [7:0] cmp289_out1;
reg [7:0] cmp289_in0;
reg [7:0] cmp289_in1;

wire [7:0] cmp290_out0;
wire [7:0] cmp290_out1;
reg [7:0] cmp290_in0;
reg [7:0] cmp290_in1;

wire [7:0] cmp291_out0;
wire [7:0] cmp291_out1;
reg [7:0] cmp291_in0;
reg [7:0] cmp291_in1;

wire [7:0] cmp292_out0;
wire [7:0] cmp292_out1;
reg [7:0] cmp292_in0;
reg [7:0] cmp292_in1;

wire [7:0] cmp293_out0;
wire [7:0] cmp293_out1;
reg [7:0] cmp293_in0;
reg [7:0] cmp293_in1;

//-------declaration layer:11----------
wire [7:0] cmp294_out0;
wire [7:0] cmp294_out1;
reg [7:0] cmp294_in0;
reg [7:0] cmp294_in1;

wire [7:0] cmp295_out0;
wire [7:0] cmp295_out1;
reg [7:0] cmp295_in0;
reg [7:0] cmp295_in1;

wire [7:0] cmp296_out0;
wire [7:0] cmp296_out1;
reg [7:0] cmp296_in0;
reg [7:0] cmp296_in1;

wire [7:0] cmp297_out0;
wire [7:0] cmp297_out1;
reg [7:0] cmp297_in0;
reg [7:0] cmp297_in1;

wire [7:0] cmp298_out0;
wire [7:0] cmp298_out1;
reg [7:0] cmp298_in0;
reg [7:0] cmp298_in1;

wire [7:0] cmp299_out0;
wire [7:0] cmp299_out1;
reg [7:0] cmp299_in0;
reg [7:0] cmp299_in1;

wire [7:0] cmp300_out0;
wire [7:0] cmp300_out1;
reg [7:0] cmp300_in0;
reg [7:0] cmp300_in1;

wire [7:0] cmp301_out0;
wire [7:0] cmp301_out1;
reg [7:0] cmp301_in0;
reg [7:0] cmp301_in1;

wire [7:0] cmp302_out0;
wire [7:0] cmp302_out1;
reg [7:0] cmp302_in0;
reg [7:0] cmp302_in1;

//-------declaration layer:12----------
wire [7:0] cmp303_out0;
wire [7:0] cmp303_out1;
reg [7:0] cmp303_in0;
reg [7:0] cmp303_in1;

wire [7:0] cmp304_out0;
wire [7:0] cmp304_out1;
reg [7:0] cmp304_in0;
reg [7:0] cmp304_in1;

wire [7:0] cmp305_out0;
wire [7:0] cmp305_out1;
reg [7:0] cmp305_in0;
reg [7:0] cmp305_in1;

wire [7:0] cmp306_out0;
wire [7:0] cmp306_out1;
reg [7:0] cmp306_in0;
reg [7:0] cmp306_in1;

wire [7:0] cmp307_out0;
wire [7:0] cmp307_out1;
reg [7:0] cmp307_in0;
reg [7:0] cmp307_in1;

wire [7:0] cmp308_out0;
wire [7:0] cmp308_out1;
reg [7:0] cmp308_in0;
reg [7:0] cmp308_in1;

wire [7:0] cmp309_out0;
wire [7:0] cmp309_out1;
reg [7:0] cmp309_in0;
reg [7:0] cmp309_in1;

wire [7:0] cmp310_out0;
wire [7:0] cmp310_out1;
reg [7:0] cmp310_in0;
reg [7:0] cmp310_in1;

wire [7:0] cmp311_out0;
wire [7:0] cmp311_out1;
reg [7:0] cmp311_in0;
reg [7:0] cmp311_in1;

wire [7:0] cmp312_out0;
wire [7:0] cmp312_out1;
reg [7:0] cmp312_in0;
reg [7:0] cmp312_in1;

wire [7:0] cmp313_out0;
wire [7:0] cmp313_out1;
reg [7:0] cmp313_in0;
reg [7:0] cmp313_in1;

wire [7:0] cmp314_out0;
wire [7:0] cmp314_out1;
reg [7:0] cmp314_in0;
reg [7:0] cmp314_in1;

wire [7:0] cmp315_out0;
wire [7:0] cmp315_out1;
reg [7:0] cmp315_in0;
reg [7:0] cmp315_in1;

wire [7:0] cmp316_out0;
wire [7:0] cmp316_out1;
reg [7:0] cmp316_in0;
reg [7:0] cmp316_in1;

wire [7:0] cmp317_out0;
wire [7:0] cmp317_out1;
reg [7:0] cmp317_in0;
reg [7:0] cmp317_in1;

wire [7:0] cmp318_out0;
wire [7:0] cmp318_out1;
reg [7:0] cmp318_in0;
reg [7:0] cmp318_in1;

wire [7:0] cmp319_out0;
wire [7:0] cmp319_out1;
reg [7:0] cmp319_in0;
reg [7:0] cmp319_in1;

wire [7:0] cmp320_out0;
wire [7:0] cmp320_out1;
reg [7:0] cmp320_in0;
reg [7:0] cmp320_in1;

wire [7:0] cmp321_out0;
wire [7:0] cmp321_out1;
reg [7:0] cmp321_in0;
reg [7:0] cmp321_in1;

wire [7:0] cmp322_out0;
wire [7:0] cmp322_out1;
reg [7:0] cmp322_in0;
reg [7:0] cmp322_in1;

wire [7:0] cmp323_out0;
wire [7:0] cmp323_out1;
reg [7:0] cmp323_in0;
reg [7:0] cmp323_in1;

wire [7:0] cmp324_out0;
wire [7:0] cmp324_out1;
reg [7:0] cmp324_in0;
reg [7:0] cmp324_in1;

wire [7:0] cmp325_out0;
wire [7:0] cmp325_out1;
reg [7:0] cmp325_in0;
reg [7:0] cmp325_in1;

wire [7:0] cmp326_out0;
wire [7:0] cmp326_out1;
reg [7:0] cmp326_in0;
reg [7:0] cmp326_in1;

wire [7:0] cmp327_out0;
wire [7:0] cmp327_out1;
reg [7:0] cmp327_in0;
reg [7:0] cmp327_in1;

//-------declaration layer:13----------
wire [7:0] cmp328_out0;
wire [7:0] cmp328_out1;
reg [7:0] cmp328_in0;
reg [7:0] cmp328_in1;

wire [7:0] cmp329_out0;
wire [7:0] cmp329_out1;
reg [7:0] cmp329_in0;
reg [7:0] cmp329_in1;

wire [7:0] cmp330_out0;
wire [7:0] cmp330_out1;
reg [7:0] cmp330_in0;
reg [7:0] cmp330_in1;

wire [7:0] cmp331_out0;
wire [7:0] cmp331_out1;
reg [7:0] cmp331_in0;
reg [7:0] cmp331_in1;

wire [7:0] cmp332_out0;
wire [7:0] cmp332_out1;
reg [7:0] cmp332_in0;
reg [7:0] cmp332_in1;

wire [7:0] cmp333_out0;
wire [7:0] cmp333_out1;
reg [7:0] cmp333_in0;
reg [7:0] cmp333_in1;

wire [7:0] cmp334_out0;
wire [7:0] cmp334_out1;
reg [7:0] cmp334_in0;
reg [7:0] cmp334_in1;

wire [7:0] cmp335_out0;
wire [7:0] cmp335_out1;
reg [7:0] cmp335_in0;
reg [7:0] cmp335_in1;

wire [7:0] cmp336_out0;
wire [7:0] cmp336_out1;
reg [7:0] cmp336_in0;
reg [7:0] cmp336_in1;

wire [7:0] cmp337_out0;
wire [7:0] cmp337_out1;
reg [7:0] cmp337_in0;
reg [7:0] cmp337_in1;

wire [7:0] cmp338_out0;
wire [7:0] cmp338_out1;
reg [7:0] cmp338_in0;
reg [7:0] cmp338_in1;

wire [7:0] cmp339_out0;
wire [7:0] cmp339_out1;
reg [7:0] cmp339_in0;
reg [7:0] cmp339_in1;

wire [7:0] cmp340_out0;
wire [7:0] cmp340_out1;
reg [7:0] cmp340_in0;
reg [7:0] cmp340_in1;

wire [7:0] cmp341_out0;
wire [7:0] cmp341_out1;
reg [7:0] cmp341_in0;
reg [7:0] cmp341_in1;

wire [7:0] cmp342_out0;
wire [7:0] cmp342_out1;
reg [7:0] cmp342_in0;
reg [7:0] cmp342_in1;

wire [7:0] cmp343_out0;
wire [7:0] cmp343_out1;
reg [7:0] cmp343_in0;
reg [7:0] cmp343_in1;

wire [7:0] cmp344_out0;
wire [7:0] cmp344_out1;
reg [7:0] cmp344_in0;
reg [7:0] cmp344_in1;

wire [7:0] cmp345_out0;
wire [7:0] cmp345_out1;
reg [7:0] cmp345_in0;
reg [7:0] cmp345_in1;

wire [7:0] cmp346_out0;
wire [7:0] cmp346_out1;
reg [7:0] cmp346_in0;
reg [7:0] cmp346_in1;

wire [7:0] cmp347_out0;
wire [7:0] cmp347_out1;
reg [7:0] cmp347_in0;
reg [7:0] cmp347_in1;

wire [7:0] cmp348_out0;
wire [7:0] cmp348_out1;
reg [7:0] cmp348_in0;
reg [7:0] cmp348_in1;

wire [7:0] cmp349_out0;
wire [7:0] cmp349_out1;
reg [7:0] cmp349_in0;
reg [7:0] cmp349_in1;

wire [7:0] cmp350_out0;
wire [7:0] cmp350_out1;
reg [7:0] cmp350_in0;
reg [7:0] cmp350_in1;

wire [7:0] cmp351_out0;
wire [7:0] cmp351_out1;
reg [7:0] cmp351_in0;
reg [7:0] cmp351_in1;

wire [7:0] cmp352_out0;
wire [7:0] cmp352_out1;
reg [7:0] cmp352_in0;
reg [7:0] cmp352_in1;

wire [7:0] cmp353_out0;
wire [7:0] cmp353_out1;
reg [7:0] cmp353_in0;
reg [7:0] cmp353_in1;

wire [7:0] cmp354_out0;
wire [7:0] cmp354_out1;
reg [7:0] cmp354_in0;
reg [7:0] cmp354_in1;

wire [7:0] cmp355_out0;
wire [7:0] cmp355_out1;
reg [7:0] cmp355_in0;
reg [7:0] cmp355_in1;

wire [7:0] cmp356_out0;
wire [7:0] cmp356_out1;
reg [7:0] cmp356_in0;
reg [7:0] cmp356_in1;

wire [7:0] cmp357_out0;
wire [7:0] cmp357_out1;
reg [7:0] cmp357_in0;
reg [7:0] cmp357_in1;

wire [7:0] cmp358_out0;
wire [7:0] cmp358_out1;
reg [7:0] cmp358_in0;
reg [7:0] cmp358_in1;

wire [7:0] cmp359_out0;
wire [7:0] cmp359_out1;
reg [7:0] cmp359_in0;
reg [7:0] cmp359_in1;

wire [7:0] cmp360_out0;
wire [7:0] cmp360_out1;
reg [7:0] cmp360_in0;
reg [7:0] cmp360_in1;

//-------declaration layer:14----------
wire [7:0] cmp361_out0;
wire [7:0] cmp361_out1;
reg [7:0] cmp361_in0;
reg [7:0] cmp361_in1;

wire [7:0] cmp362_out0;
wire [7:0] cmp362_out1;
reg [7:0] cmp362_in0;
reg [7:0] cmp362_in1;

wire [7:0] cmp363_out0;
wire [7:0] cmp363_out1;
reg [7:0] cmp363_in0;
reg [7:0] cmp363_in1;

wire [7:0] cmp364_out0;
wire [7:0] cmp364_out1;
reg [7:0] cmp364_in0;
reg [7:0] cmp364_in1;

wire [7:0] cmp365_out0;
wire [7:0] cmp365_out1;
reg [7:0] cmp365_in0;
reg [7:0] cmp365_in1;

wire [7:0] cmp366_out0;
wire [7:0] cmp366_out1;
reg [7:0] cmp366_in0;
reg [7:0] cmp366_in1;

wire [7:0] cmp367_out0;
wire [7:0] cmp367_out1;
reg [7:0] cmp367_in0;
reg [7:0] cmp367_in1;

wire [7:0] cmp368_out0;
wire [7:0] cmp368_out1;
reg [7:0] cmp368_in0;
reg [7:0] cmp368_in1;

wire [7:0] cmp369_out0;
wire [7:0] cmp369_out1;
reg [7:0] cmp369_in0;
reg [7:0] cmp369_in1;

wire [7:0] cmp370_out0;
wire [7:0] cmp370_out1;
reg [7:0] cmp370_in0;
reg [7:0] cmp370_in1;

wire [7:0] cmp371_out0;
wire [7:0] cmp371_out1;
reg [7:0] cmp371_in0;
reg [7:0] cmp371_in1;

wire [7:0] cmp372_out0;
wire [7:0] cmp372_out1;
reg [7:0] cmp372_in0;
reg [7:0] cmp372_in1;

wire [7:0] cmp373_out0;
wire [7:0] cmp373_out1;
reg [7:0] cmp373_in0;
reg [7:0] cmp373_in1;

wire [7:0] cmp374_out0;
wire [7:0] cmp374_out1;
reg [7:0] cmp374_in0;
reg [7:0] cmp374_in1;

wire [7:0] cmp375_out0;
wire [7:0] cmp375_out1;
reg [7:0] cmp375_in0;
reg [7:0] cmp375_in1;

wire [7:0] cmp376_out0;
wire [7:0] cmp376_out1;
reg [7:0] cmp376_in0;
reg [7:0] cmp376_in1;

wire [7:0] cmp377_out0;
wire [7:0] cmp377_out1;
reg [7:0] cmp377_in0;
reg [7:0] cmp377_in1;

wire [7:0] cmp378_out0;
wire [7:0] cmp378_out1;
reg [7:0] cmp378_in0;
reg [7:0] cmp378_in1;

wire [7:0] cmp379_out0;
wire [7:0] cmp379_out1;
reg [7:0] cmp379_in0;
reg [7:0] cmp379_in1;

wire [7:0] cmp380_out0;
wire [7:0] cmp380_out1;
reg [7:0] cmp380_in0;
reg [7:0] cmp380_in1;

wire [7:0] cmp381_out0;
wire [7:0] cmp381_out1;
reg [7:0] cmp381_in0;
reg [7:0] cmp381_in1;

wire [7:0] cmp382_out0;
wire [7:0] cmp382_out1;
reg [7:0] cmp382_in0;
reg [7:0] cmp382_in1;

wire [7:0] cmp383_out0;
wire [7:0] cmp383_out1;
reg [7:0] cmp383_in0;
reg [7:0] cmp383_in1;

wire [7:0] cmp384_out0;
wire [7:0] cmp384_out1;
reg [7:0] cmp384_in0;
reg [7:0] cmp384_in1;

wire [7:0] cmp385_out0;
wire [7:0] cmp385_out1;
reg [7:0] cmp385_in0;
reg [7:0] cmp385_in1;

wire [7:0] cmp386_out0;
wire [7:0] cmp386_out1;
reg [7:0] cmp386_in0;
reg [7:0] cmp386_in1;

wire [7:0] cmp387_out0;
wire [7:0] cmp387_out1;
reg [7:0] cmp387_in0;
reg [7:0] cmp387_in1;

wire [7:0] cmp388_out0;
wire [7:0] cmp388_out1;
reg [7:0] cmp388_in0;
reg [7:0] cmp388_in1;

wire [7:0] cmp389_out0;
wire [7:0] cmp389_out1;
reg [7:0] cmp389_in0;
reg [7:0] cmp389_in1;

wire [7:0] cmp390_out0;
wire [7:0] cmp390_out1;
reg [7:0] cmp390_in0;
reg [7:0] cmp390_in1;

wire [7:0] cmp391_out0;
wire [7:0] cmp391_out1;
reg [7:0] cmp391_in0;
reg [7:0] cmp391_in1;

wire [7:0] cmp392_out0;
wire [7:0] cmp392_out1;
reg [7:0] cmp392_in0;
reg [7:0] cmp392_in1;

wire [7:0] cmp393_out0;
wire [7:0] cmp393_out1;
reg [7:0] cmp393_in0;
reg [7:0] cmp393_in1;

wire [7:0] cmp394_out0;
wire [7:0] cmp394_out1;
reg [7:0] cmp394_in0;
reg [7:0] cmp394_in1;

wire [7:0] cmp395_out0;
wire [7:0] cmp395_out1;
reg [7:0] cmp395_in0;
reg [7:0] cmp395_in1;

wire [7:0] cmp396_out0;
wire [7:0] cmp396_out1;
reg [7:0] cmp396_in0;
reg [7:0] cmp396_in1;

wire [7:0] cmp397_out0;
wire [7:0] cmp397_out1;
reg [7:0] cmp397_in0;
reg [7:0] cmp397_in1;

wire [7:0] cmp398_out0;
wire [7:0] cmp398_out1;
reg [7:0] cmp398_in0;
reg [7:0] cmp398_in1;

wire [7:0] cmp399_out0;
wire [7:0] cmp399_out1;
reg [7:0] cmp399_in0;
reg [7:0] cmp399_in1;

//-------declaration layer:15----------
wire [7:0] cmp400_out0;
wire [7:0] cmp400_out1;
reg [7:0] cmp400_in0;
reg [7:0] cmp400_in1;

wire [7:0] cmp401_out0;
wire [7:0] cmp401_out1;
reg [7:0] cmp401_in0;
reg [7:0] cmp401_in1;

wire [7:0] cmp402_out0;
wire [7:0] cmp402_out1;
reg [7:0] cmp402_in0;
reg [7:0] cmp402_in1;

wire [7:0] cmp403_out0;
wire [7:0] cmp403_out1;
reg [7:0] cmp403_in0;
reg [7:0] cmp403_in1;

wire [7:0] cmp404_out0;
wire [7:0] cmp404_out1;
reg [7:0] cmp404_in0;
reg [7:0] cmp404_in1;

wire [7:0] cmp405_out0;
wire [7:0] cmp405_out1;
reg [7:0] cmp405_in0;
reg [7:0] cmp405_in1;

wire [7:0] cmp406_out0;
wire [7:0] cmp406_out1;
reg [7:0] cmp406_in0;
reg [7:0] cmp406_in1;

wire [7:0] cmp407_out0;
wire [7:0] cmp407_out1;
reg [7:0] cmp407_in0;
reg [7:0] cmp407_in1;

wire [7:0] cmp408_out0;
wire [7:0] cmp408_out1;
reg [7:0] cmp408_in0;
reg [7:0] cmp408_in1;

wire [7:0] cmp409_out0;
wire [7:0] cmp409_out1;
reg [7:0] cmp409_in0;
reg [7:0] cmp409_in1;

wire [7:0] cmp410_out0;
wire [7:0] cmp410_out1;
reg [7:0] cmp410_in0;
reg [7:0] cmp410_in1;

wire [7:0] cmp411_out0;
wire [7:0] cmp411_out1;
reg [7:0] cmp411_in0;
reg [7:0] cmp411_in1;

wire [7:0] cmp412_out0;
wire [7:0] cmp412_out1;
reg [7:0] cmp412_in0;
reg [7:0] cmp412_in1;

wire [7:0] cmp413_out0;
wire [7:0] cmp413_out1;
reg [7:0] cmp413_in0;
reg [7:0] cmp413_in1;

wire [7:0] cmp414_out0;
wire [7:0] cmp414_out1;
reg [7:0] cmp414_in0;
reg [7:0] cmp414_in1;

wire [7:0] cmp415_out0;
wire [7:0] cmp415_out1;
reg [7:0] cmp415_in0;
reg [7:0] cmp415_in1;

wire [7:0] cmp416_out0;
wire [7:0] cmp416_out1;
reg [7:0] cmp416_in0;
reg [7:0] cmp416_in1;

wire [7:0] cmp417_out0;
wire [7:0] cmp417_out1;
reg [7:0] cmp417_in0;
reg [7:0] cmp417_in1;

wire [7:0] cmp418_out0;
wire [7:0] cmp418_out1;
reg [7:0] cmp418_in0;
reg [7:0] cmp418_in1;

wire [7:0] cmp419_out0;
wire [7:0] cmp419_out1;
reg [7:0] cmp419_in0;
reg [7:0] cmp419_in1;

wire [7:0] cmp420_out0;
wire [7:0] cmp420_out1;
reg [7:0] cmp420_in0;
reg [7:0] cmp420_in1;

wire [7:0] cmp421_out0;
wire [7:0] cmp421_out1;
reg [7:0] cmp421_in0;
reg [7:0] cmp421_in1;

wire [7:0] cmp422_out0;
wire [7:0] cmp422_out1;
reg [7:0] cmp422_in0;
reg [7:0] cmp422_in1;

wire [7:0] cmp423_out0;
wire [7:0] cmp423_out1;
reg [7:0] cmp423_in0;
reg [7:0] cmp423_in1;

wire [7:0] cmp424_out0;
wire [7:0] cmp424_out1;
reg [7:0] cmp424_in0;
reg [7:0] cmp424_in1;

wire [7:0] cmp425_out0;
wire [7:0] cmp425_out1;
reg [7:0] cmp425_in0;
reg [7:0] cmp425_in1;

wire [7:0] cmp426_out0;
wire [7:0] cmp426_out1;
reg [7:0] cmp426_in0;
reg [7:0] cmp426_in1;

wire [7:0] cmp427_out0;
wire [7:0] cmp427_out1;
reg [7:0] cmp427_in0;
reg [7:0] cmp427_in1;

wire [7:0] cmp428_out0;
wire [7:0] cmp428_out1;
reg [7:0] cmp428_in0;
reg [7:0] cmp428_in1;

wire [7:0] cmp429_out0;
wire [7:0] cmp429_out1;
reg [7:0] cmp429_in0;
reg [7:0] cmp429_in1;

wire [7:0] cmp430_out0;
wire [7:0] cmp430_out1;
reg [7:0] cmp430_in0;
reg [7:0] cmp430_in1;

wire [7:0] cmp431_out0;
wire [7:0] cmp431_out1;
reg [7:0] cmp431_in0;
reg [7:0] cmp431_in1;

wire [7:0] cmp432_out0;
wire [7:0] cmp432_out1;
reg [7:0] cmp432_in0;
reg [7:0] cmp432_in1;

wire [7:0] cmp433_out0;
wire [7:0] cmp433_out1;
reg [7:0] cmp433_in0;
reg [7:0] cmp433_in1;

wire [7:0] cmp434_out0;
wire [7:0] cmp434_out1;
reg [7:0] cmp434_in0;
reg [7:0] cmp434_in1;

wire [7:0] cmp435_out0;
wire [7:0] cmp435_out1;
reg [7:0] cmp435_in0;
reg [7:0] cmp435_in1;

wire [7:0] cmp436_out0;
wire [7:0] cmp436_out1;
reg [7:0] cmp436_in0;
reg [7:0] cmp436_in1;

wire [7:0] cmp437_out0;
wire [7:0] cmp437_out1;
reg [7:0] cmp437_in0;
reg [7:0] cmp437_in1;

//-------declaration layer:16----------
wire [7:0] cmp438_out0;
wire [7:0] cmp438_out1;
reg [7:0] cmp438_in0;
reg [7:0] cmp438_in1;

wire [7:0] cmp439_out0;
wire [7:0] cmp439_out1;
reg [7:0] cmp439_in0;
reg [7:0] cmp439_in1;

wire [7:0] cmp440_out0;
wire [7:0] cmp440_out1;
reg [7:0] cmp440_in0;
reg [7:0] cmp440_in1;

wire [7:0] cmp441_out0;
wire [7:0] cmp441_out1;
reg [7:0] cmp441_in0;
reg [7:0] cmp441_in1;

wire [7:0] cmp442_out0;
wire [7:0] cmp442_out1;
reg [7:0] cmp442_in0;
reg [7:0] cmp442_in1;

wire [7:0] cmp443_out0;
wire [7:0] cmp443_out1;
reg [7:0] cmp443_in0;
reg [7:0] cmp443_in1;

wire [7:0] cmp444_out0;
wire [7:0] cmp444_out1;
reg [7:0] cmp444_in0;
reg [7:0] cmp444_in1;

wire [7:0] cmp445_out0;
wire [7:0] cmp445_out1;
reg [7:0] cmp445_in0;
reg [7:0] cmp445_in1;

wire [7:0] cmp446_out0;
wire [7:0] cmp446_out1;
reg [7:0] cmp446_in0;
reg [7:0] cmp446_in1;

//-------declaration layer:17----------
wire [7:0] cmp447_out0;
wire [7:0] cmp447_out1;
reg [7:0] cmp447_in0;
reg [7:0] cmp447_in1;

wire [7:0] cmp448_out0;
wire [7:0] cmp448_out1;
reg [7:0] cmp448_in0;
reg [7:0] cmp448_in1;

wire [7:0] cmp449_out0;
wire [7:0] cmp449_out1;
reg [7:0] cmp449_in0;
reg [7:0] cmp449_in1;

wire [7:0] cmp450_out0;
wire [7:0] cmp450_out1;
reg [7:0] cmp450_in0;
reg [7:0] cmp450_in1;

wire [7:0] cmp451_out0;
wire [7:0] cmp451_out1;
reg [7:0] cmp451_in0;
reg [7:0] cmp451_in1;

wire [7:0] cmp452_out0;
wire [7:0] cmp452_out1;
reg [7:0] cmp452_in0;
reg [7:0] cmp452_in1;

wire [7:0] cmp453_out0;
wire [7:0] cmp453_out1;
reg [7:0] cmp453_in0;
reg [7:0] cmp453_in1;

wire [7:0] cmp454_out0;
wire [7:0] cmp454_out1;
reg [7:0] cmp454_in0;
reg [7:0] cmp454_in1;

wire [7:0] cmp455_out0;
wire [7:0] cmp455_out1;
reg [7:0] cmp455_in0;
reg [7:0] cmp455_in1;

wire [7:0] cmp456_out0;
wire [7:0] cmp456_out1;
reg [7:0] cmp456_in0;
reg [7:0] cmp456_in1;

wire [7:0] cmp457_out0;
wire [7:0] cmp457_out1;
reg [7:0] cmp457_in0;
reg [7:0] cmp457_in1;

wire [7:0] cmp458_out0;
wire [7:0] cmp458_out1;
reg [7:0] cmp458_in0;
reg [7:0] cmp458_in1;

wire [7:0] cmp459_out0;
wire [7:0] cmp459_out1;
reg [7:0] cmp459_in0;
reg [7:0] cmp459_in1;

wire [7:0] cmp460_out0;
wire [7:0] cmp460_out1;
reg [7:0] cmp460_in0;
reg [7:0] cmp460_in1;

wire [7:0] cmp461_out0;
wire [7:0] cmp461_out1;
reg [7:0] cmp461_in0;
reg [7:0] cmp461_in1;

wire [7:0] cmp462_out0;
wire [7:0] cmp462_out1;
reg [7:0] cmp462_in0;
reg [7:0] cmp462_in1;

wire [7:0] cmp463_out0;
wire [7:0] cmp463_out1;
reg [7:0] cmp463_in0;
reg [7:0] cmp463_in1;

wire [7:0] cmp464_out0;
wire [7:0] cmp464_out1;
reg [7:0] cmp464_in0;
reg [7:0] cmp464_in1;

wire [7:0] cmp465_out0;
wire [7:0] cmp465_out1;
reg [7:0] cmp465_in0;
reg [7:0] cmp465_in1;

wire [7:0] cmp466_out0;
wire [7:0] cmp466_out1;
reg [7:0] cmp466_in0;
reg [7:0] cmp466_in1;

wire [7:0] cmp467_out0;
wire [7:0] cmp467_out1;
reg [7:0] cmp467_in0;
reg [7:0] cmp467_in1;

wire [7:0] cmp468_out0;
wire [7:0] cmp468_out1;
reg [7:0] cmp468_in0;
reg [7:0] cmp468_in1;

wire [7:0] cmp469_out0;
wire [7:0] cmp469_out1;
reg [7:0] cmp469_in0;
reg [7:0] cmp469_in1;

wire [7:0] cmp470_out0;
wire [7:0] cmp470_out1;
reg [7:0] cmp470_in0;
reg [7:0] cmp470_in1;

wire [7:0] cmp471_out0;
wire [7:0] cmp471_out1;
reg [7:0] cmp471_in0;
reg [7:0] cmp471_in1;

//-------declaration layer:18----------
wire [7:0] cmp472_out0;
wire [7:0] cmp472_out1;
reg [7:0] cmp472_in0;
reg [7:0] cmp472_in1;

wire [7:0] cmp473_out0;
wire [7:0] cmp473_out1;
reg [7:0] cmp473_in0;
reg [7:0] cmp473_in1;

wire [7:0] cmp474_out0;
wire [7:0] cmp474_out1;
reg [7:0] cmp474_in0;
reg [7:0] cmp474_in1;

wire [7:0] cmp475_out0;
wire [7:0] cmp475_out1;
reg [7:0] cmp475_in0;
reg [7:0] cmp475_in1;

wire [7:0] cmp476_out0;
wire [7:0] cmp476_out1;
reg [7:0] cmp476_in0;
reg [7:0] cmp476_in1;

wire [7:0] cmp477_out0;
wire [7:0] cmp477_out1;
reg [7:0] cmp477_in0;
reg [7:0] cmp477_in1;

wire [7:0] cmp478_out0;
wire [7:0] cmp478_out1;
reg [7:0] cmp478_in0;
reg [7:0] cmp478_in1;

wire [7:0] cmp479_out0;
wire [7:0] cmp479_out1;
reg [7:0] cmp479_in0;
reg [7:0] cmp479_in1;

wire [7:0] cmp480_out0;
wire [7:0] cmp480_out1;
reg [7:0] cmp480_in0;
reg [7:0] cmp480_in1;

wire [7:0] cmp481_out0;
wire [7:0] cmp481_out1;
reg [7:0] cmp481_in0;
reg [7:0] cmp481_in1;

wire [7:0] cmp482_out0;
wire [7:0] cmp482_out1;
reg [7:0] cmp482_in0;
reg [7:0] cmp482_in1;

wire [7:0] cmp483_out0;
wire [7:0] cmp483_out1;
reg [7:0] cmp483_in0;
reg [7:0] cmp483_in1;

wire [7:0] cmp484_out0;
wire [7:0] cmp484_out1;
reg [7:0] cmp484_in0;
reg [7:0] cmp484_in1;

wire [7:0] cmp485_out0;
wire [7:0] cmp485_out1;
reg [7:0] cmp485_in0;
reg [7:0] cmp485_in1;

wire [7:0] cmp486_out0;
wire [7:0] cmp486_out1;
reg [7:0] cmp486_in0;
reg [7:0] cmp486_in1;

wire [7:0] cmp487_out0;
wire [7:0] cmp487_out1;
reg [7:0] cmp487_in0;
reg [7:0] cmp487_in1;

wire [7:0] cmp488_out0;
wire [7:0] cmp488_out1;
reg [7:0] cmp488_in0;
reg [7:0] cmp488_in1;

wire [7:0] cmp489_out0;
wire [7:0] cmp489_out1;
reg [7:0] cmp489_in0;
reg [7:0] cmp489_in1;

wire [7:0] cmp490_out0;
wire [7:0] cmp490_out1;
reg [7:0] cmp490_in0;
reg [7:0] cmp490_in1;

wire [7:0] cmp491_out0;
wire [7:0] cmp491_out1;
reg [7:0] cmp491_in0;
reg [7:0] cmp491_in1;

wire [7:0] cmp492_out0;
wire [7:0] cmp492_out1;
reg [7:0] cmp492_in0;
reg [7:0] cmp492_in1;

wire [7:0] cmp493_out0;
wire [7:0] cmp493_out1;
reg [7:0] cmp493_in0;
reg [7:0] cmp493_in1;

wire [7:0] cmp494_out0;
wire [7:0] cmp494_out1;
reg [7:0] cmp494_in0;
reg [7:0] cmp494_in1;

wire [7:0] cmp495_out0;
wire [7:0] cmp495_out1;
reg [7:0] cmp495_in0;
reg [7:0] cmp495_in1;

wire [7:0] cmp496_out0;
wire [7:0] cmp496_out1;
reg [7:0] cmp496_in0;
reg [7:0] cmp496_in1;

wire [7:0] cmp497_out0;
wire [7:0] cmp497_out1;
reg [7:0] cmp497_in0;
reg [7:0] cmp497_in1;

wire [7:0] cmp498_out0;
wire [7:0] cmp498_out1;
reg [7:0] cmp498_in0;
reg [7:0] cmp498_in1;

wire [7:0] cmp499_out0;
wire [7:0] cmp499_out1;
reg [7:0] cmp499_in0;
reg [7:0] cmp499_in1;

wire [7:0] cmp500_out0;
wire [7:0] cmp500_out1;
reg [7:0] cmp500_in0;
reg [7:0] cmp500_in1;

wire [7:0] cmp501_out0;
wire [7:0] cmp501_out1;
reg [7:0] cmp501_in0;
reg [7:0] cmp501_in1;

wire [7:0] cmp502_out0;
wire [7:0] cmp502_out1;
reg [7:0] cmp502_in0;
reg [7:0] cmp502_in1;

wire [7:0] cmp503_out0;
wire [7:0] cmp503_out1;
reg [7:0] cmp503_in0;
reg [7:0] cmp503_in1;

wire [7:0] cmp504_out0;
wire [7:0] cmp504_out1;
reg [7:0] cmp504_in0;
reg [7:0] cmp504_in1;

//-------declaration layer:19----------
wire [7:0] cmp505_out0;
wire [7:0] cmp505_out1;
reg [7:0] cmp505_in0;
reg [7:0] cmp505_in1;

wire [7:0] cmp506_out0;
wire [7:0] cmp506_out1;
reg [7:0] cmp506_in0;
reg [7:0] cmp506_in1;

wire [7:0] cmp507_out0;
wire [7:0] cmp507_out1;
reg [7:0] cmp507_in0;
reg [7:0] cmp507_in1;

wire [7:0] cmp508_out0;
wire [7:0] cmp508_out1;
reg [7:0] cmp508_in0;
reg [7:0] cmp508_in1;

wire [7:0] cmp509_out0;
wire [7:0] cmp509_out1;
reg [7:0] cmp509_in0;
reg [7:0] cmp509_in1;

wire [7:0] cmp510_out0;
wire [7:0] cmp510_out1;
reg [7:0] cmp510_in0;
reg [7:0] cmp510_in1;

wire [7:0] cmp511_out0;
wire [7:0] cmp511_out1;
reg [7:0] cmp511_in0;
reg [7:0] cmp511_in1;

wire [7:0] cmp512_out0;
wire [7:0] cmp512_out1;
reg [7:0] cmp512_in0;
reg [7:0] cmp512_in1;

wire [7:0] cmp513_out0;
wire [7:0] cmp513_out1;
reg [7:0] cmp513_in0;
reg [7:0] cmp513_in1;

wire [7:0] cmp514_out0;
wire [7:0] cmp514_out1;
reg [7:0] cmp514_in0;
reg [7:0] cmp514_in1;

wire [7:0] cmp515_out0;
wire [7:0] cmp515_out1;
reg [7:0] cmp515_in0;
reg [7:0] cmp515_in1;

wire [7:0] cmp516_out0;
wire [7:0] cmp516_out1;
reg [7:0] cmp516_in0;
reg [7:0] cmp516_in1;

wire [7:0] cmp517_out0;
wire [7:0] cmp517_out1;
reg [7:0] cmp517_in0;
reg [7:0] cmp517_in1;

wire [7:0] cmp518_out0;
wire [7:0] cmp518_out1;
reg [7:0] cmp518_in0;
reg [7:0] cmp518_in1;

wire [7:0] cmp519_out0;
wire [7:0] cmp519_out1;
reg [7:0] cmp519_in0;
reg [7:0] cmp519_in1;

wire [7:0] cmp520_out0;
wire [7:0] cmp520_out1;
reg [7:0] cmp520_in0;
reg [7:0] cmp520_in1;

wire [7:0] cmp521_out0;
wire [7:0] cmp521_out1;
reg [7:0] cmp521_in0;
reg [7:0] cmp521_in1;

wire [7:0] cmp522_out0;
wire [7:0] cmp522_out1;
reg [7:0] cmp522_in0;
reg [7:0] cmp522_in1;

wire [7:0] cmp523_out0;
wire [7:0] cmp523_out1;
reg [7:0] cmp523_in0;
reg [7:0] cmp523_in1;

wire [7:0] cmp524_out0;
wire [7:0] cmp524_out1;
reg [7:0] cmp524_in0;
reg [7:0] cmp524_in1;

wire [7:0] cmp525_out0;
wire [7:0] cmp525_out1;
reg [7:0] cmp525_in0;
reg [7:0] cmp525_in1;

wire [7:0] cmp526_out0;
wire [7:0] cmp526_out1;
reg [7:0] cmp526_in0;
reg [7:0] cmp526_in1;

wire [7:0] cmp527_out0;
wire [7:0] cmp527_out1;
reg [7:0] cmp527_in0;
reg [7:0] cmp527_in1;

wire [7:0] cmp528_out0;
wire [7:0] cmp528_out1;
reg [7:0] cmp528_in0;
reg [7:0] cmp528_in1;

wire [7:0] cmp529_out0;
wire [7:0] cmp529_out1;
reg [7:0] cmp529_in0;
reg [7:0] cmp529_in1;

wire [7:0] cmp530_out0;
wire [7:0] cmp530_out1;
reg [7:0] cmp530_in0;
reg [7:0] cmp530_in1;

wire [7:0] cmp531_out0;
wire [7:0] cmp531_out1;
reg [7:0] cmp531_in0;
reg [7:0] cmp531_in1;

wire [7:0] cmp532_out0;
wire [7:0] cmp532_out1;
reg [7:0] cmp532_in0;
reg [7:0] cmp532_in1;

wire [7:0] cmp533_out0;
wire [7:0] cmp533_out1;
reg [7:0] cmp533_in0;
reg [7:0] cmp533_in1;

wire [7:0] cmp534_out0;
wire [7:0] cmp534_out1;
reg [7:0] cmp534_in0;
reg [7:0] cmp534_in1;

wire [7:0] cmp535_out0;
wire [7:0] cmp535_out1;
reg [7:0] cmp535_in0;
reg [7:0] cmp535_in1;

wire [7:0] cmp536_out0;
wire [7:0] cmp536_out1;
reg [7:0] cmp536_in0;
reg [7:0] cmp536_in1;

wire [7:0] cmp537_out0;
wire [7:0] cmp537_out1;
reg [7:0] cmp537_in0;
reg [7:0] cmp537_in1;

wire [7:0] cmp538_out0;
wire [7:0] cmp538_out1;
reg [7:0] cmp538_in0;
reg [7:0] cmp538_in1;

wire [7:0] cmp539_out0;
wire [7:0] cmp539_out1;
reg [7:0] cmp539_in0;
reg [7:0] cmp539_in1;

wire [7:0] cmp540_out0;
wire [7:0] cmp540_out1;
reg [7:0] cmp540_in0;
reg [7:0] cmp540_in1;

wire [7:0] cmp541_out0;
wire [7:0] cmp541_out1;
reg [7:0] cmp541_in0;
reg [7:0] cmp541_in1;

//-------declaration layer:20----------
wire [7:0] cmp542_out0;
wire [7:0] cmp542_out1;
reg [7:0] cmp542_in0;
reg [7:0] cmp542_in1;

wire [7:0] cmp543_out0;
wire [7:0] cmp543_out1;
reg [7:0] cmp543_in0;
reg [7:0] cmp543_in1;

wire [7:0] cmp544_out0;
wire [7:0] cmp544_out1;
reg [7:0] cmp544_in0;
reg [7:0] cmp544_in1;

wire [7:0] cmp545_out0;
wire [7:0] cmp545_out1;
reg [7:0] cmp545_in0;
reg [7:0] cmp545_in1;

wire [7:0] cmp546_out0;
wire [7:0] cmp546_out1;
reg [7:0] cmp546_in0;
reg [7:0] cmp546_in1;

wire [7:0] cmp547_out0;
wire [7:0] cmp547_out1;
reg [7:0] cmp547_in0;
reg [7:0] cmp547_in1;

wire [7:0] cmp548_out0;
wire [7:0] cmp548_out1;
reg [7:0] cmp548_in0;
reg [7:0] cmp548_in1;

wire [7:0] cmp549_out0;
wire [7:0] cmp549_out1;
reg [7:0] cmp549_in0;
reg [7:0] cmp549_in1;

wire [7:0] cmp550_out0;
wire [7:0] cmp550_out1;
reg [7:0] cmp550_in0;
reg [7:0] cmp550_in1;

wire [7:0] cmp551_out0;
wire [7:0] cmp551_out1;
reg [7:0] cmp551_in0;
reg [7:0] cmp551_in1;

wire [7:0] cmp552_out0;
wire [7:0] cmp552_out1;
reg [7:0] cmp552_in0;
reg [7:0] cmp552_in1;

wire [7:0] cmp553_out0;
wire [7:0] cmp553_out1;
reg [7:0] cmp553_in0;
reg [7:0] cmp553_in1;

wire [7:0] cmp554_out0;
wire [7:0] cmp554_out1;
reg [7:0] cmp554_in0;
reg [7:0] cmp554_in1;

wire [7:0] cmp555_out0;
wire [7:0] cmp555_out1;
reg [7:0] cmp555_in0;
reg [7:0] cmp555_in1;

wire [7:0] cmp556_out0;
wire [7:0] cmp556_out1;
reg [7:0] cmp556_in0;
reg [7:0] cmp556_in1;

wire [7:0] cmp557_out0;
wire [7:0] cmp557_out1;
reg [7:0] cmp557_in0;
reg [7:0] cmp557_in1;

wire [7:0] cmp558_out0;
wire [7:0] cmp558_out1;
reg [7:0] cmp558_in0;
reg [7:0] cmp558_in1;

wire [7:0] cmp559_out0;
wire [7:0] cmp559_out1;
reg [7:0] cmp559_in0;
reg [7:0] cmp559_in1;

wire [7:0] cmp560_out0;
wire [7:0] cmp560_out1;
reg [7:0] cmp560_in0;
reg [7:0] cmp560_in1;

wire [7:0] cmp561_out0;
wire [7:0] cmp561_out1;
reg [7:0] cmp561_in0;
reg [7:0] cmp561_in1;

wire [7:0] cmp562_out0;
wire [7:0] cmp562_out1;
reg [7:0] cmp562_in0;
reg [7:0] cmp562_in1;

wire [7:0] cmp563_out0;
wire [7:0] cmp563_out1;
reg [7:0] cmp563_in0;
reg [7:0] cmp563_in1;

wire [7:0] cmp564_out0;
wire [7:0] cmp564_out1;
reg [7:0] cmp564_in0;
reg [7:0] cmp564_in1;

wire [7:0] cmp565_out0;
wire [7:0] cmp565_out1;
reg [7:0] cmp565_in0;
reg [7:0] cmp565_in1;

wire [7:0] cmp566_out0;
wire [7:0] cmp566_out1;
reg [7:0] cmp566_in0;
reg [7:0] cmp566_in1;

wire [7:0] cmp567_out0;
wire [7:0] cmp567_out1;
reg [7:0] cmp567_in0;
reg [7:0] cmp567_in1;

wire [7:0] cmp568_out0;
wire [7:0] cmp568_out1;
reg [7:0] cmp568_in0;
reg [7:0] cmp568_in1;

wire [7:0] cmp569_out0;
wire [7:0] cmp569_out1;
reg [7:0] cmp569_in0;
reg [7:0] cmp569_in1;

wire [7:0] cmp570_out0;
wire [7:0] cmp570_out1;
reg [7:0] cmp570_in0;
reg [7:0] cmp570_in1;

wire [7:0] cmp571_out0;
wire [7:0] cmp571_out1;
reg [7:0] cmp571_in0;
reg [7:0] cmp571_in1;

wire [7:0] cmp572_out0;
wire [7:0] cmp572_out1;
reg [7:0] cmp572_in0;
reg [7:0] cmp572_in1;

wire [7:0] cmp573_out0;
wire [7:0] cmp573_out1;
reg [7:0] cmp573_in0;
reg [7:0] cmp573_in1;

wire [7:0] cmp574_out0;
wire [7:0] cmp574_out1;
reg [7:0] cmp574_in0;
reg [7:0] cmp574_in1;

wire [7:0] cmp575_out0;
wire [7:0] cmp575_out1;
reg [7:0] cmp575_in0;
reg [7:0] cmp575_in1;

wire [7:0] cmp576_out0;
wire [7:0] cmp576_out1;
reg [7:0] cmp576_in0;
reg [7:0] cmp576_in1;

wire [7:0] cmp577_out0;
wire [7:0] cmp577_out1;
reg [7:0] cmp577_in0;
reg [7:0] cmp577_in1;

wire [7:0] cmp578_out0;
wire [7:0] cmp578_out1;
reg [7:0] cmp578_in0;
reg [7:0] cmp578_in1;

wire [7:0] cmp579_out0;
wire [7:0] cmp579_out1;
reg [7:0] cmp579_in0;
reg [7:0] cmp579_in1;

wire [7:0] cmp580_out0;
wire [7:0] cmp580_out1;
reg [7:0] cmp580_in0;
reg [7:0] cmp580_in1;

wire [7:0] cmp581_out0;
wire [7:0] cmp581_out1;
reg [7:0] cmp581_in0;
reg [7:0] cmp581_in1;

//-------declaration layer:21----------
wire [7:0] cmp582_out0;
wire [7:0] cmp582_out1;
reg [7:0] cmp582_in0;
reg [7:0] cmp582_in1;

wire [7:0] cmp583_out0;
wire [7:0] cmp583_out1;
reg [7:0] cmp583_in0;
reg [7:0] cmp583_in1;

wire [7:0] cmp584_out0;
wire [7:0] cmp584_out1;
reg [7:0] cmp584_in0;
reg [7:0] cmp584_in1;

wire [7:0] cmp585_out0;
wire [7:0] cmp585_out1;
reg [7:0] cmp585_in0;
reg [7:0] cmp585_in1;

wire [7:0] cmp586_out0;
wire [7:0] cmp586_out1;
reg [7:0] cmp586_in0;
reg [7:0] cmp586_in1;

wire [7:0] cmp587_out0;
wire [7:0] cmp587_out1;
reg [7:0] cmp587_in0;
reg [7:0] cmp587_in1;

wire [7:0] cmp588_out0;
wire [7:0] cmp588_out1;
reg [7:0] cmp588_in0;
reg [7:0] cmp588_in1;

wire [7:0] cmp589_out0;
wire [7:0] cmp589_out1;
reg [7:0] cmp589_in0;
reg [7:0] cmp589_in1;

wire [7:0] cmp590_out0;
wire [7:0] cmp590_out1;
reg [7:0] cmp590_in0;
reg [7:0] cmp590_in1;

wire [7:0] cmp591_out0;
wire [7:0] cmp591_out1;
reg [7:0] cmp591_in0;
reg [7:0] cmp591_in1;

wire [7:0] cmp592_out0;
wire [7:0] cmp592_out1;
reg [7:0] cmp592_in0;
reg [7:0] cmp592_in1;

wire [7:0] cmp593_out0;
wire [7:0] cmp593_out1;
reg [7:0] cmp593_in0;
reg [7:0] cmp593_in1;

wire [7:0] cmp594_out0;
wire [7:0] cmp594_out1;
reg [7:0] cmp594_in0;
reg [7:0] cmp594_in1;

wire [7:0] cmp595_out0;
wire [7:0] cmp595_out1;
reg [7:0] cmp595_in0;
reg [7:0] cmp595_in1;

wire [7:0] cmp596_out0;
wire [7:0] cmp596_out1;
reg [7:0] cmp596_in0;
reg [7:0] cmp596_in1;

wire [7:0] cmp597_out0;
wire [7:0] cmp597_out1;
reg [7:0] cmp597_in0;
reg [7:0] cmp597_in1;

wire [7:0] cmp598_out0;
wire [7:0] cmp598_out1;
reg [7:0] cmp598_in0;
reg [7:0] cmp598_in1;

wire [7:0] cmp599_out0;
wire [7:0] cmp599_out1;
reg [7:0] cmp599_in0;
reg [7:0] cmp599_in1;

wire [7:0] cmp600_out0;
wire [7:0] cmp600_out1;
reg [7:0] cmp600_in0;
reg [7:0] cmp600_in1;

wire [7:0] cmp601_out0;
wire [7:0] cmp601_out1;
reg [7:0] cmp601_in0;
reg [7:0] cmp601_in1;

wire [7:0] cmp602_out0;
wire [7:0] cmp602_out1;
reg [7:0] cmp602_in0;
reg [7:0] cmp602_in1;

wire [7:0] cmp603_out0;
wire [7:0] cmp603_out1;
reg [7:0] cmp603_in0;
reg [7:0] cmp603_in1;

wire [7:0] cmp604_out0;
wire [7:0] cmp604_out1;
reg [7:0] cmp604_in0;
reg [7:0] cmp604_in1;

wire [7:0] cmp605_out0;
wire [7:0] cmp605_out1;
reg [7:0] cmp605_in0;
reg [7:0] cmp605_in1;

wire [7:0] cmp606_out0;
wire [7:0] cmp606_out1;
reg [7:0] cmp606_in0;
reg [7:0] cmp606_in1;

wire [7:0] cmp607_out0;
wire [7:0] cmp607_out1;
reg [7:0] cmp607_in0;
reg [7:0] cmp607_in1;

wire [7:0] cmp608_out0;
wire [7:0] cmp608_out1;
reg [7:0] cmp608_in0;
reg [7:0] cmp608_in1;

wire [7:0] cmp609_out0;
wire [7:0] cmp609_out1;
reg [7:0] cmp609_in0;
reg [7:0] cmp609_in1;

wire [7:0] cmp610_out0;
wire [7:0] cmp610_out1;
reg [7:0] cmp610_in0;
reg [7:0] cmp610_in1;

wire [7:0] cmp611_out0;
wire [7:0] cmp611_out1;
reg [7:0] cmp611_in0;
reg [7:0] cmp611_in1;

wire [7:0] cmp612_out0;
wire [7:0] cmp612_out1;
reg [7:0] cmp612_in0;
reg [7:0] cmp612_in1;

wire [7:0] cmp613_out0;
wire [7:0] cmp613_out1;
reg [7:0] cmp613_in0;
reg [7:0] cmp613_in1;

wire [7:0] cmp614_out0;
wire [7:0] cmp614_out1;
reg [7:0] cmp614_in0;
reg [7:0] cmp614_in1;

wire [7:0] cmp615_out0;
wire [7:0] cmp615_out1;
reg [7:0] cmp615_in0;
reg [7:0] cmp615_in1;

wire [7:0] cmp616_out0;
wire [7:0] cmp616_out1;
reg [7:0] cmp616_in0;
reg [7:0] cmp616_in1;

wire [7:0] cmp617_out0;
wire [7:0] cmp617_out1;
reg [7:0] cmp617_in0;
reg [7:0] cmp617_in1;

wire [7:0] cmp618_out0;
wire [7:0] cmp618_out1;
reg [7:0] cmp618_in0;
reg [7:0] cmp618_in1;

wire [7:0] cmp619_out0;
wire [7:0] cmp619_out1;
reg [7:0] cmp619_in0;
reg [7:0] cmp619_in1;

wire [7:0] cmp620_out0;
wire [7:0] cmp620_out1;
reg [7:0] cmp620_in0;
reg [7:0] cmp620_in1;

//-------declaration layer:22----------
wire [7:0] cmp621_out0;
wire [7:0] cmp621_out1;
reg [7:0] cmp621_in0;
reg [7:0] cmp621_in1;

wire [7:0] cmp622_out0;
wire [7:0] cmp622_out1;
reg [7:0] cmp622_in0;
reg [7:0] cmp622_in1;

wire [7:0] cmp623_out0;
wire [7:0] cmp623_out1;
reg [7:0] cmp623_in0;
reg [7:0] cmp623_in1;

wire [7:0] cmp624_out0;
wire [7:0] cmp624_out1;
reg [7:0] cmp624_in0;
reg [7:0] cmp624_in1;

wire [7:0] cmp625_out0;
wire [7:0] cmp625_out1;
reg [7:0] cmp625_in0;
reg [7:0] cmp625_in1;

wire [7:0] cmp626_out0;
wire [7:0] cmp626_out1;
reg [7:0] cmp626_in0;
reg [7:0] cmp626_in1;

wire [7:0] cmp627_out0;
wire [7:0] cmp627_out1;
reg [7:0] cmp627_in0;
reg [7:0] cmp627_in1;

wire [7:0] cmp628_out0;
wire [7:0] cmp628_out1;
reg [7:0] cmp628_in0;
reg [7:0] cmp628_in1;

wire [7:0] cmp629_out0;
wire [7:0] cmp629_out1;
reg [7:0] cmp629_in0;
reg [7:0] cmp629_in1;

//-------declaration layer:23----------
wire [7:0] cmp630_out0;
wire [7:0] cmp630_out1;
reg [7:0] cmp630_in0;
reg [7:0] cmp630_in1;

wire [7:0] cmp631_out0;
wire [7:0] cmp631_out1;
reg [7:0] cmp631_in0;
reg [7:0] cmp631_in1;

wire [7:0] cmp632_out0;
wire [7:0] cmp632_out1;
reg [7:0] cmp632_in0;
reg [7:0] cmp632_in1;

wire [7:0] cmp633_out0;
wire [7:0] cmp633_out1;
reg [7:0] cmp633_in0;
reg [7:0] cmp633_in1;

wire [7:0] cmp634_out0;
wire [7:0] cmp634_out1;
reg [7:0] cmp634_in0;
reg [7:0] cmp634_in1;

wire [7:0] cmp635_out0;
wire [7:0] cmp635_out1;
reg [7:0] cmp635_in0;
reg [7:0] cmp635_in1;

wire [7:0] cmp636_out0;
wire [7:0] cmp636_out1;
reg [7:0] cmp636_in0;
reg [7:0] cmp636_in1;

wire [7:0] cmp637_out0;
wire [7:0] cmp637_out1;
reg [7:0] cmp637_in0;
reg [7:0] cmp637_in1;

wire [7:0] cmp638_out0;
wire [7:0] cmp638_out1;
reg [7:0] cmp638_in0;
reg [7:0] cmp638_in1;

wire [7:0] cmp639_out0;
wire [7:0] cmp639_out1;
reg [7:0] cmp639_in0;
reg [7:0] cmp639_in1;

wire [7:0] cmp640_out0;
wire [7:0] cmp640_out1;
reg [7:0] cmp640_in0;
reg [7:0] cmp640_in1;

wire [7:0] cmp641_out0;
wire [7:0] cmp641_out1;
reg [7:0] cmp641_in0;
reg [7:0] cmp641_in1;

wire [7:0] cmp642_out0;
wire [7:0] cmp642_out1;
reg [7:0] cmp642_in0;
reg [7:0] cmp642_in1;

wire [7:0] cmp643_out0;
wire [7:0] cmp643_out1;
reg [7:0] cmp643_in0;
reg [7:0] cmp643_in1;

wire [7:0] cmp644_out0;
wire [7:0] cmp644_out1;
reg [7:0] cmp644_in0;
reg [7:0] cmp644_in1;

wire [7:0] cmp645_out0;
wire [7:0] cmp645_out1;
reg [7:0] cmp645_in0;
reg [7:0] cmp645_in1;

//-------declaration layer:24----------
wire [7:0] cmp646_out0;
wire [7:0] cmp646_out1;
reg [7:0] cmp646_in0;
reg [7:0] cmp646_in1;

wire [7:0] cmp647_out0;
wire [7:0] cmp647_out1;
reg [7:0] cmp647_in0;
reg [7:0] cmp647_in1;

wire [7:0] cmp648_out0;
wire [7:0] cmp648_out1;
reg [7:0] cmp648_in0;
reg [7:0] cmp648_in1;

wire [7:0] cmp649_out0;
wire [7:0] cmp649_out1;
reg [7:0] cmp649_in0;
reg [7:0] cmp649_in1;

wire [7:0] cmp650_out0;
wire [7:0] cmp650_out1;
reg [7:0] cmp650_in0;
reg [7:0] cmp650_in1;

wire [7:0] cmp651_out0;
wire [7:0] cmp651_out1;
reg [7:0] cmp651_in0;
reg [7:0] cmp651_in1;

wire [7:0] cmp652_out0;
wire [7:0] cmp652_out1;
reg [7:0] cmp652_in0;
reg [7:0] cmp652_in1;

wire [7:0] cmp653_out0;
wire [7:0] cmp653_out1;
reg [7:0] cmp653_in0;
reg [7:0] cmp653_in1;

//-------declaration layer:25----------
wire [7:0] cmp654_out0;
wire [7:0] cmp654_out1;
reg [7:0] cmp654_in0;
reg [7:0] cmp654_in1;

wire [7:0] cmp655_out0;
wire [7:0] cmp655_out1;
reg [7:0] cmp655_in0;
reg [7:0] cmp655_in1;

wire [7:0] cmp656_out0;
wire [7:0] cmp656_out1;
reg [7:0] cmp656_in0;
reg [7:0] cmp656_in1;

wire [7:0] cmp657_out0;
wire [7:0] cmp657_out1;
reg [7:0] cmp657_in0;
reg [7:0] cmp657_in1;

//-------declaration layer:26----------
wire [7:0] cmp658_out0;
wire [7:0] cmp658_out1;
reg [7:0] cmp658_in0;
reg [7:0] cmp658_in1;

wire [7:0] cmp659_out0;
wire [7:0] cmp659_out1;
reg [7:0] cmp659_in0;
reg [7:0] cmp659_in1;

//-------declaration layer:27----------
wire [7:0] cmp660_out0;
wire [7:0] cmp660_out1;
reg [7:0] cmp660_in0;
reg [7:0] cmp660_in1;

//-------Temp Register----------
reg [7:0] r0_17_tmp;
reg [7:0] r0_18_tmp;
reg [7:0] r0_19_tmp;
reg [7:0] r0_20_tmp;
reg [7:0] r0_21_tmp;
reg [7:0] r0_22_tmp;
reg [7:0] r0_23_tmp;
reg [7:0] r0_24_tmp;
reg [7:0] r0_25_tmp;
reg [7:0] r0_26_tmp;
reg [7:0] r0_27_tmp;
reg [7:0] r0_28_tmp;
reg [7:0] r0_29_tmp;
reg [7:0] r0_30_tmp;
reg [7:0] r0_31_tmp;
reg [7:0] r0_32_tmp;
reg [7:0] r0_33_tmp;
reg [7:0] r0_34_tmp;
reg [7:0] r0_35_tmp;
reg [7:0] r0_36_tmp;
reg [7:0] r0_37_tmp;
reg [7:0] r0_38_tmp;
reg [7:0] r0_39_tmp;
reg [7:0] r0_40_tmp;
reg [7:0] r0_41_tmp;
reg [7:0] r0_42_tmp;
reg [7:0] r0_43_tmp;
reg [7:0] r0_44_tmp;
reg [7:0] r0_45_tmp;
reg [7:0] r0_46_tmp;
reg [7:0] r0_47_tmp;
reg [7:0] r0_48_tmp;
reg [7:0] r0_49_tmp;
reg [7:0] r0_50_tmp;
reg [7:0] r0_51_tmp;
reg [7:0] r0_52_tmp;
reg [7:0] r0_53_tmp;
reg [7:0] r0_54_tmp;
reg [7:0] r0_55_tmp;
reg [7:0] r0_56_tmp;
reg [7:0] r0_57_tmp;
reg [7:0] r0_58_tmp;
reg [7:0] r0_59_tmp;
reg [7:0] r0_60_tmp;
reg [7:0] r0_61_tmp;
reg [7:0] r0_62_tmp;
reg [7:0] r0_63_tmp;
reg [7:0] r1_64_tmp;
reg [7:0] r1_65_tmp;
reg [7:0] r1_66_tmp;
reg [7:0] r1_67_tmp;
reg [7:0] r1_68_tmp;
reg [7:0] r1_69_tmp;
reg [7:0] r1_70_tmp;
reg [7:0] r1_71_tmp;
reg [7:0] r1_72_tmp;
reg [7:0] r1_73_tmp;
reg [7:0] r1_74_tmp;
reg [7:0] r1_75_tmp;
reg [7:0] r1_76_tmp;
reg [7:0] r1_77_tmp;
reg [7:0] r1_78_tmp;
reg [7:0] r1_79_tmp;
reg [7:0] r1_80_tmp;
reg [7:0] r2_49_tmp;
reg [7:0] r2_50_tmp;
reg [7:0] r2_51_tmp;
reg [7:0] r2_52_tmp;
reg [7:0] r2_53_tmp;
reg [7:0] r2_54_tmp;
reg [7:0] r2_55_tmp;
reg [7:0] r2_56_tmp;
reg [7:0] r2_57_tmp;
reg [7:0] r2_58_tmp;
reg [7:0] r2_59_tmp;
reg [7:0] r2_60_tmp;
reg [7:0] r2_61_tmp;
reg [7:0] r2_62_tmp;
reg [7:0] r2_63_tmp;
reg [7:0] r3_0_tmp;
reg [7:0] r3_1_tmp;
reg [7:0] r3_2_tmp;
reg [7:0] r3_3_tmp;
reg [7:0] r3_4_tmp;
reg [7:0] r3_5_tmp;
reg [7:0] r3_6_tmp;
reg [7:0] r3_7_tmp;
reg [7:0] r3_8_tmp;
reg [7:0] r3_9_tmp;
reg [7:0] r3_10_tmp;
reg [7:0] r3_11_tmp;
reg [7:0] r3_12_tmp;
reg [7:0] r3_13_tmp;
reg [7:0] r3_14_tmp;
reg [7:0] r3_15_tmp;
reg [7:0] r3_16_tmp;
reg [7:0] r3_17_tmp;
reg [7:0] r3_18_tmp;
reg [7:0] r3_19_tmp;
reg [7:0] r3_20_tmp;
reg [7:0] r3_21_tmp;
reg [7:0] r3_22_tmp;
reg [7:0] r3_23_tmp;
reg [7:0] r3_24_tmp;
reg [7:0] r3_25_tmp;
reg [7:0] r3_26_tmp;
reg [7:0] r3_27_tmp;
reg [7:0] r3_28_tmp;
reg [7:0] r3_29_tmp;
reg [7:0] r3_30_tmp;
reg [7:0] r3_31_tmp;
reg [7:0] r3_65_tmp;
reg [7:0] r3_66_tmp;
reg [7:0] r3_67_tmp;
reg [7:0] r3_68_tmp;
reg [7:0] r3_69_tmp;
reg [7:0] r3_70_tmp;
reg [7:0] r3_71_tmp;
reg [7:0] r3_72_tmp;
reg [7:0] r3_73_tmp;
reg [7:0] r3_74_tmp;
reg [7:0] r3_75_tmp;
reg [7:0] r3_76_tmp;
reg [7:0] r3_77_tmp;
reg [7:0] r3_78_tmp;
reg [7:0] r3_79_tmp;
reg [7:0] r4_0_tmp;
reg [7:0] r4_1_tmp;
reg [7:0] r4_2_tmp;
reg [7:0] r4_3_tmp;
reg [7:0] r4_4_tmp;
reg [7:0] r4_5_tmp;
reg [7:0] r4_6_tmp;
reg [7:0] r4_7_tmp;
reg [7:0] r4_8_tmp;
reg [7:0] r4_9_tmp;
reg [7:0] r4_10_tmp;
reg [7:0] r4_11_tmp;
reg [7:0] r4_12_tmp;
reg [7:0] r4_13_tmp;
reg [7:0] r4_14_tmp;
reg [7:0] r4_15_tmp;
reg [7:0] r4_32_tmp;
reg [7:0] r4_33_tmp;
reg [7:0] r4_34_tmp;
reg [7:0] r4_35_tmp;
reg [7:0] r4_36_tmp;
reg [7:0] r4_37_tmp;
reg [7:0] r4_38_tmp;
reg [7:0] r4_39_tmp;
reg [7:0] r4_40_tmp;
reg [7:0] r4_41_tmp;
reg [7:0] r4_42_tmp;
reg [7:0] r4_43_tmp;
reg [7:0] r4_44_tmp;
reg [7:0] r4_45_tmp;
reg [7:0] r4_46_tmp;
reg [7:0] r4_47_tmp;
reg [7:0] r4_48_tmp;
reg [7:0] r4_49_tmp;
reg [7:0] r4_50_tmp;
reg [7:0] r4_51_tmp;
reg [7:0] r4_52_tmp;
reg [7:0] r4_53_tmp;
reg [7:0] r4_54_tmp;
reg [7:0] r4_55_tmp;
reg [7:0] r4_56_tmp;
reg [7:0] r4_57_tmp;
reg [7:0] r4_58_tmp;
reg [7:0] r4_59_tmp;
reg [7:0] r4_60_tmp;
reg [7:0] r4_61_tmp;
reg [7:0] r4_62_tmp;
reg [7:0] r4_63_tmp;
reg [7:0] r4_80_tmp;
reg [7:0] r5_80_tmp;
reg [7:0] r6_0_tmp;
reg [7:0] r6_1_tmp;
reg [7:0] r6_2_tmp;
reg [7:0] r6_3_tmp;
reg [7:0] r6_4_tmp;
reg [7:0] r6_5_tmp;
reg [7:0] r6_6_tmp;
reg [7:0] r6_7_tmp;
reg [7:0] r6_8_tmp;
reg [7:0] r6_9_tmp;
reg [7:0] r6_10_tmp;
reg [7:0] r6_11_tmp;
reg [7:0] r6_12_tmp;
reg [7:0] r6_13_tmp;
reg [7:0] r6_14_tmp;
reg [7:0] r6_15_tmp;
reg [7:0] r6_80_tmp;
reg [7:0] r7_0_tmp;
reg [7:0] r7_1_tmp;
reg [7:0] r7_2_tmp;
reg [7:0] r7_3_tmp;
reg [7:0] r7_4_tmp;
reg [7:0] r7_5_tmp;
reg [7:0] r7_6_tmp;
reg [7:0] r7_7_tmp;
reg [7:0] r7_16_tmp;
reg [7:0] r7_17_tmp;
reg [7:0] r7_18_tmp;
reg [7:0] r7_19_tmp;
reg [7:0] r7_20_tmp;
reg [7:0] r7_21_tmp;
reg [7:0] r7_22_tmp;
reg [7:0] r7_23_tmp;
reg [7:0] r7_25_tmp;
reg [7:0] r7_26_tmp;
reg [7:0] r7_27_tmp;
reg [7:0] r7_28_tmp;
reg [7:0] r7_29_tmp;
reg [7:0] r7_30_tmp;
reg [7:0] r7_31_tmp;
reg [7:0] r7_32_tmp;
reg [7:0] r7_33_tmp;
reg [7:0] r7_34_tmp;
reg [7:0] r7_35_tmp;
reg [7:0] r7_36_tmp;
reg [7:0] r7_37_tmp;
reg [7:0] r7_38_tmp;
reg [7:0] r7_39_tmp;
reg [7:0] r7_40_tmp;
reg [7:0] r7_41_tmp;
reg [7:0] r7_42_tmp;
reg [7:0] r7_43_tmp;
reg [7:0] r7_44_tmp;
reg [7:0] r7_45_tmp;
reg [7:0] r7_46_tmp;
reg [7:0] r7_47_tmp;
reg [7:0] r7_48_tmp;
reg [7:0] r7_49_tmp;
reg [7:0] r7_50_tmp;
reg [7:0] r7_51_tmp;
reg [7:0] r7_52_tmp;
reg [7:0] r7_53_tmp;
reg [7:0] r7_54_tmp;
reg [7:0] r7_55_tmp;
reg [7:0] r7_56_tmp;
reg [7:0] r7_57_tmp;
reg [7:0] r7_58_tmp;
reg [7:0] r7_59_tmp;
reg [7:0] r7_60_tmp;
reg [7:0] r7_61_tmp;
reg [7:0] r7_62_tmp;
reg [7:0] r7_63_tmp;
reg [7:0] r7_72_tmp;
reg [7:0] r7_73_tmp;
reg [7:0] r7_74_tmp;
reg [7:0] r7_75_tmp;
reg [7:0] r7_76_tmp;
reg [7:0] r7_77_tmp;
reg [7:0] r7_78_tmp;
reg [7:0] r7_79_tmp;
reg [7:0] r8_0_tmp;
reg [7:0] r8_1_tmp;
reg [7:0] r8_2_tmp;
reg [7:0] r8_3_tmp;
reg [7:0] r8_4_tmp;
reg [7:0] r8_5_tmp;
reg [7:0] r8_6_tmp;
reg [7:0] r8_7_tmp;
reg [7:0] r8_16_tmp;
reg [7:0] r8_17_tmp;
reg [7:0] r8_18_tmp;
reg [7:0] r8_19_tmp;
reg [7:0] r8_20_tmp;
reg [7:0] r8_21_tmp;
reg [7:0] r8_22_tmp;
reg [7:0] r8_23_tmp;
reg [7:0] r8_57_tmp;
reg [7:0] r8_58_tmp;
reg [7:0] r8_59_tmp;
reg [7:0] r8_60_tmp;
reg [7:0] r8_61_tmp;
reg [7:0] r8_62_tmp;
reg [7:0] r8_63_tmp;
reg [7:0] r8_72_tmp;
reg [7:0] r8_73_tmp;
reg [7:0] r8_74_tmp;
reg [7:0] r8_75_tmp;
reg [7:0] r8_76_tmp;
reg [7:0] r8_77_tmp;
reg [7:0] r8_78_tmp;
reg [7:0] r8_79_tmp;
reg [7:0] r9_73_tmp;
reg [7:0] r9_74_tmp;
reg [7:0] r9_75_tmp;
reg [7:0] r9_76_tmp;
reg [7:0] r9_77_tmp;
reg [7:0] r9_78_tmp;
reg [7:0] r9_79_tmp;
reg [7:0] r10_0_tmp;
reg [7:0] r10_1_tmp;
reg [7:0] r10_2_tmp;
reg [7:0] r10_3_tmp;
reg [7:0] r10_4_tmp;
reg [7:0] r10_5_tmp;
reg [7:0] r10_6_tmp;
reg [7:0] r10_7_tmp;
reg [7:0] r10_80_tmp;
reg [7:0] r11_0_tmp;
reg [7:0] r11_1_tmp;
reg [7:0] r11_2_tmp;
reg [7:0] r11_3_tmp;
reg [7:0] r11_8_tmp;
reg [7:0] r11_9_tmp;
reg [7:0] r11_10_tmp;
reg [7:0] r11_11_tmp;
reg [7:0] r11_16_tmp;
reg [7:0] r11_17_tmp;
reg [7:0] r11_18_tmp;
reg [7:0] r11_19_tmp;
reg [7:0] r11_21_tmp;
reg [7:0] r11_22_tmp;
reg [7:0] r11_23_tmp;
reg [7:0] r11_24_tmp;
reg [7:0] r11_25_tmp;
reg [7:0] r11_26_tmp;
reg [7:0] r11_27_tmp;
reg [7:0] r11_28_tmp;
reg [7:0] r11_29_tmp;
reg [7:0] r11_30_tmp;
reg [7:0] r11_31_tmp;
reg [7:0] r11_32_tmp;
reg [7:0] r11_33_tmp;
reg [7:0] r11_34_tmp;
reg [7:0] r11_35_tmp;
reg [7:0] r11_36_tmp;
reg [7:0] r11_37_tmp;
reg [7:0] r11_38_tmp;
reg [7:0] r11_39_tmp;
reg [7:0] r11_40_tmp;
reg [7:0] r11_41_tmp;
reg [7:0] r11_42_tmp;
reg [7:0] r11_43_tmp;
reg [7:0] r11_44_tmp;
reg [7:0] r11_45_tmp;
reg [7:0] r11_46_tmp;
reg [7:0] r11_47_tmp;
reg [7:0] r11_48_tmp;
reg [7:0] r11_49_tmp;
reg [7:0] r11_50_tmp;
reg [7:0] r11_51_tmp;
reg [7:0] r11_52_tmp;
reg [7:0] r11_53_tmp;
reg [7:0] r11_54_tmp;
reg [7:0] r11_55_tmp;
reg [7:0] r11_56_tmp;
reg [7:0] r11_57_tmp;
reg [7:0] r11_58_tmp;
reg [7:0] r11_59_tmp;
reg [7:0] r11_60_tmp;
reg [7:0] r11_61_tmp;
reg [7:0] r11_62_tmp;
reg [7:0] r11_63_tmp;
reg [7:0] r11_68_tmp;
reg [7:0] r11_69_tmp;
reg [7:0] r11_70_tmp;
reg [7:0] r11_71_tmp;
reg [7:0] r11_76_tmp;
reg [7:0] r11_77_tmp;
reg [7:0] r11_78_tmp;
reg [7:0] r11_79_tmp;
reg [7:0] r12_0_tmp;
reg [7:0] r12_1_tmp;
reg [7:0] r12_2_tmp;
reg [7:0] r12_3_tmp;
reg [7:0] r12_8_tmp;
reg [7:0] r12_9_tmp;
reg [7:0] r12_10_tmp;
reg [7:0] r12_11_tmp;
reg [7:0] r12_16_tmp;
reg [7:0] r12_17_tmp;
reg [7:0] r12_18_tmp;
reg [7:0] r12_19_tmp;
reg [7:0] r12_24_tmp;
reg [7:0] r12_25_tmp;
reg [7:0] r12_26_tmp;
reg [7:0] r12_27_tmp;
reg [7:0] r12_53_tmp;
reg [7:0] r12_54_tmp;
reg [7:0] r12_55_tmp;
reg [7:0] r12_60_tmp;
reg [7:0] r12_61_tmp;
reg [7:0] r12_62_tmp;
reg [7:0] r12_63_tmp;
reg [7:0] r12_68_tmp;
reg [7:0] r12_69_tmp;
reg [7:0] r12_70_tmp;
reg [7:0] r12_71_tmp;
reg [7:0] r12_76_tmp;
reg [7:0] r12_77_tmp;
reg [7:0] r12_78_tmp;
reg [7:0] r12_79_tmp;
reg [7:0] r13_0_tmp;
reg [7:0] r13_1_tmp;
reg [7:0] r13_2_tmp;
reg [7:0] r13_3_tmp;
reg [7:0] r13_8_tmp;
reg [7:0] r13_9_tmp;
reg [7:0] r13_10_tmp;
reg [7:0] r13_11_tmp;
reg [7:0] r13_69_tmp;
reg [7:0] r13_70_tmp;
reg [7:0] r13_71_tmp;
reg [7:0] r13_76_tmp;
reg [7:0] r13_77_tmp;
reg [7:0] r13_78_tmp;
reg [7:0] r13_79_tmp;
reg [7:0] r14_77_tmp;
reg [7:0] r14_78_tmp;
reg [7:0] r14_79_tmp;
reg [7:0] r15_0_tmp;
reg [7:0] r15_1_tmp;
reg [7:0] r15_2_tmp;
reg [7:0] r15_3_tmp;
reg [7:0] r15_80_tmp;
reg [7:0] r16_0_tmp;
reg [7:0] r16_1_tmp;
reg [7:0] r16_4_tmp;
reg [7:0] r16_5_tmp;
reg [7:0] r16_8_tmp;
reg [7:0] r16_9_tmp;
reg [7:0] r16_12_tmp;
reg [7:0] r16_13_tmp;
reg [7:0] r16_16_tmp;
reg [7:0] r16_17_tmp;
reg [7:0] r16_19_tmp;
reg [7:0] r16_20_tmp;
reg [7:0] r16_21_tmp;
reg [7:0] r16_22_tmp;
reg [7:0] r16_23_tmp;
reg [7:0] r16_24_tmp;
reg [7:0] r16_25_tmp;
reg [7:0] r16_26_tmp;
reg [7:0] r16_27_tmp;
reg [7:0] r16_28_tmp;
reg [7:0] r16_29_tmp;
reg [7:0] r16_30_tmp;
reg [7:0] r16_31_tmp;
reg [7:0] r16_32_tmp;
reg [7:0] r16_33_tmp;
reg [7:0] r16_34_tmp;
reg [7:0] r16_35_tmp;
reg [7:0] r16_36_tmp;
reg [7:0] r16_37_tmp;
reg [7:0] r16_38_tmp;
reg [7:0] r16_39_tmp;
reg [7:0] r16_40_tmp;
reg [7:0] r16_41_tmp;
reg [7:0] r16_42_tmp;
reg [7:0] r16_43_tmp;
reg [7:0] r16_44_tmp;
reg [7:0] r16_45_tmp;
reg [7:0] r16_46_tmp;
reg [7:0] r16_47_tmp;
reg [7:0] r16_48_tmp;
reg [7:0] r16_49_tmp;
reg [7:0] r16_50_tmp;
reg [7:0] r16_51_tmp;
reg [7:0] r16_52_tmp;
reg [7:0] r16_53_tmp;
reg [7:0] r16_54_tmp;
reg [7:0] r16_55_tmp;
reg [7:0] r16_56_tmp;
reg [7:0] r16_57_tmp;
reg [7:0] r16_58_tmp;
reg [7:0] r16_59_tmp;
reg [7:0] r16_60_tmp;
reg [7:0] r16_61_tmp;
reg [7:0] r16_62_tmp;
reg [7:0] r16_63_tmp;
reg [7:0] r16_66_tmp;
reg [7:0] r16_67_tmp;
reg [7:0] r16_70_tmp;
reg [7:0] r16_71_tmp;
reg [7:0] r16_74_tmp;
reg [7:0] r16_75_tmp;
reg [7:0] r16_78_tmp;
reg [7:0] r16_79_tmp;
reg [7:0] r17_0_tmp;
reg [7:0] r17_1_tmp;
reg [7:0] r17_4_tmp;
reg [7:0] r17_5_tmp;
reg [7:0] r17_8_tmp;
reg [7:0] r17_9_tmp;
reg [7:0] r17_12_tmp;
reg [7:0] r17_13_tmp;
reg [7:0] r17_16_tmp;
reg [7:0] r17_17_tmp;
reg [7:0] r17_20_tmp;
reg [7:0] r17_21_tmp;
reg [7:0] r17_24_tmp;
reg [7:0] r17_25_tmp;
reg [7:0] r17_28_tmp;
reg [7:0] r17_29_tmp;
reg [7:0] r17_51_tmp;
reg [7:0] r17_54_tmp;
reg [7:0] r17_55_tmp;
reg [7:0] r17_58_tmp;
reg [7:0] r17_59_tmp;
reg [7:0] r17_62_tmp;
reg [7:0] r17_63_tmp;
reg [7:0] r17_66_tmp;
reg [7:0] r17_67_tmp;
reg [7:0] r17_70_tmp;
reg [7:0] r17_71_tmp;
reg [7:0] r17_74_tmp;
reg [7:0] r17_75_tmp;
reg [7:0] r17_78_tmp;
reg [7:0] r17_79_tmp;
reg [7:0] r18_0_tmp;
reg [7:0] r18_1_tmp;
reg [7:0] r18_4_tmp;
reg [7:0] r18_5_tmp;
reg [7:0] r18_8_tmp;
reg [7:0] r18_9_tmp;
reg [7:0] r18_12_tmp;
reg [7:0] r18_13_tmp;
reg [7:0] r18_67_tmp;
reg [7:0] r18_70_tmp;
reg [7:0] r18_71_tmp;
reg [7:0] r18_74_tmp;
reg [7:0] r18_75_tmp;
reg [7:0] r18_78_tmp;
reg [7:0] r18_79_tmp;
reg [7:0] r19_0_tmp;
reg [7:0] r19_1_tmp;
reg [7:0] r19_4_tmp;
reg [7:0] r19_5_tmp;
reg [7:0] r19_75_tmp;
reg [7:0] r19_78_tmp;
reg [7:0] r19_79_tmp;
reg [7:0] r20_79_tmp;
reg [7:0] r21_0_tmp;
reg [7:0] r21_1_tmp;
reg [7:0] r21_80_tmp;
reg [7:0] r22_0_tmp;
reg [7:0] r22_2_tmp;
reg [7:0] r22_4_tmp;
reg [7:0] r22_6_tmp;
reg [7:0] r22_8_tmp;
reg [7:0] r22_10_tmp;
reg [7:0] r22_12_tmp;
reg [7:0] r22_14_tmp;
reg [7:0] r22_16_tmp;
reg [7:0] r22_18_tmp;
reg [7:0] r22_19_tmp;
reg [7:0] r22_20_tmp;
reg [7:0] r22_21_tmp;
reg [7:0] r22_22_tmp;
reg [7:0] r22_23_tmp;
reg [7:0] r22_24_tmp;
reg [7:0] r22_25_tmp;
reg [7:0] r22_26_tmp;
reg [7:0] r22_27_tmp;
reg [7:0] r22_28_tmp;
reg [7:0] r22_29_tmp;
reg [7:0] r22_30_tmp;
reg [7:0] r22_31_tmp;
reg [7:0] r22_32_tmp;
reg [7:0] r22_33_tmp;
reg [7:0] r22_34_tmp;
reg [7:0] r22_35_tmp;
reg [7:0] r22_36_tmp;
reg [7:0] r22_37_tmp;
reg [7:0] r22_38_tmp;
reg [7:0] r22_39_tmp;
reg [7:0] r22_40_tmp;
reg [7:0] r22_41_tmp;
reg [7:0] r22_42_tmp;
reg [7:0] r22_43_tmp;
reg [7:0] r22_44_tmp;
reg [7:0] r22_45_tmp;
reg [7:0] r22_46_tmp;
reg [7:0] r22_47_tmp;
reg [7:0] r22_48_tmp;
reg [7:0] r22_49_tmp;
reg [7:0] r22_50_tmp;
reg [7:0] r22_51_tmp;
reg [7:0] r22_52_tmp;
reg [7:0] r22_53_tmp;
reg [7:0] r22_54_tmp;
reg [7:0] r22_55_tmp;
reg [7:0] r22_56_tmp;
reg [7:0] r22_57_tmp;
reg [7:0] r22_58_tmp;
reg [7:0] r22_59_tmp;
reg [7:0] r22_60_tmp;
reg [7:0] r22_61_tmp;
reg [7:0] r22_62_tmp;
reg [7:0] r22_63_tmp;
reg [7:0] r22_65_tmp;
reg [7:0] r22_67_tmp;
reg [7:0] r22_69_tmp;
reg [7:0] r22_71_tmp;
reg [7:0] r22_73_tmp;
reg [7:0] r22_75_tmp;
reg [7:0] r22_77_tmp;
reg [7:0] r22_79_tmp;
reg [7:0] r23_0_tmp;
reg [7:0] r23_1_tmp;
reg [7:0] r23_2_tmp;
reg [7:0] r23_3_tmp;
reg [7:0] r23_4_tmp;
reg [7:0] r23_5_tmp;
reg [7:0] r23_6_tmp;
reg [7:0] r23_7_tmp;
reg [7:0] r23_8_tmp;
reg [7:0] r23_10_tmp;
reg [7:0] r23_12_tmp;
reg [7:0] r23_14_tmp;
reg [7:0] r23_16_tmp;
reg [7:0] r23_18_tmp;
reg [7:0] r23_20_tmp;
reg [7:0] r23_22_tmp;
reg [7:0] r23_24_tmp;
reg [7:0] r23_26_tmp;
reg [7:0] r23_28_tmp;
reg [7:0] r23_30_tmp;
reg [7:0] r23_32_tmp;
reg [7:0] r23_34_tmp;
reg [7:0] r23_36_tmp;
reg [7:0] r23_38_tmp;
reg [7:0] r23_41_tmp;
reg [7:0] r23_43_tmp;
reg [7:0] r23_45_tmp;
reg [7:0] r23_47_tmp;
reg [7:0] r23_49_tmp;
reg [7:0] r23_51_tmp;
reg [7:0] r23_53_tmp;
reg [7:0] r23_55_tmp;
reg [7:0] r23_57_tmp;
reg [7:0] r23_59_tmp;
reg [7:0] r23_61_tmp;
reg [7:0] r23_63_tmp;
reg [7:0] r23_65_tmp;
reg [7:0] r23_67_tmp;
reg [7:0] r23_69_tmp;
reg [7:0] r23_71_tmp;
reg [7:0] r23_72_tmp;
reg [7:0] r23_73_tmp;
reg [7:0] r23_74_tmp;
reg [7:0] r23_75_tmp;
reg [7:0] r23_76_tmp;
reg [7:0] r23_77_tmp;
reg [7:0] r23_78_tmp;
reg [7:0] r23_79_tmp;
reg [7:0] r23_80_tmp;
reg [7:0] r24_0_tmp;
reg [7:0] r24_1_tmp;
reg [7:0] r24_2_tmp;
reg [7:0] r24_3_tmp;
reg [7:0] r24_4_tmp;
reg [7:0] r24_5_tmp;
reg [7:0] r24_6_tmp;
reg [7:0] r24_7_tmp;
reg [7:0] r24_8_tmp;
reg [7:0] r24_9_tmp;
reg [7:0] r24_10_tmp;
reg [7:0] r24_11_tmp;
reg [7:0] r24_12_tmp;
reg [7:0] r24_13_tmp;
reg [7:0] r24_14_tmp;
reg [7:0] r24_15_tmp;
reg [7:0] r24_16_tmp;
reg [7:0] r24_17_tmp;
reg [7:0] r24_18_tmp;
reg [7:0] r24_19_tmp;
reg [7:0] r24_20_tmp;
reg [7:0] r24_21_tmp;
reg [7:0] r24_22_tmp;
reg [7:0] r24_23_tmp;
reg [7:0] r24_24_tmp;
reg [7:0] r24_26_tmp;
reg [7:0] r24_28_tmp;
reg [7:0] r24_30_tmp;
reg [7:0] r24_32_tmp;
reg [7:0] r24_34_tmp;
reg [7:0] r24_36_tmp;
reg [7:0] r24_38_tmp;
reg [7:0] r24_41_tmp;
reg [7:0] r24_43_tmp;
reg [7:0] r24_45_tmp;
reg [7:0] r24_47_tmp;
reg [7:0] r24_49_tmp;
reg [7:0] r24_51_tmp;
reg [7:0] r24_53_tmp;
reg [7:0] r24_55_tmp;
reg [7:0] r24_56_tmp;
reg [7:0] r24_57_tmp;
reg [7:0] r24_58_tmp;
reg [7:0] r24_59_tmp;
reg [7:0] r24_60_tmp;
reg [7:0] r24_61_tmp;
reg [7:0] r24_62_tmp;
reg [7:0] r24_63_tmp;
reg [7:0] r24_64_tmp;
reg [7:0] r24_65_tmp;
reg [7:0] r24_66_tmp;
reg [7:0] r24_67_tmp;
reg [7:0] r24_68_tmp;
reg [7:0] r24_69_tmp;
reg [7:0] r24_70_tmp;
reg [7:0] r24_71_tmp;
reg [7:0] r24_72_tmp;
reg [7:0] r24_73_tmp;
reg [7:0] r24_74_tmp;
reg [7:0] r24_75_tmp;
reg [7:0] r24_76_tmp;
reg [7:0] r24_77_tmp;
reg [7:0] r24_78_tmp;
reg [7:0] r24_79_tmp;
reg [7:0] r24_80_tmp;
reg [7:0] r25_0_tmp;
reg [7:0] r25_1_tmp;
reg [7:0] r25_2_tmp;
reg [7:0] r25_3_tmp;
reg [7:0] r25_4_tmp;
reg [7:0] r25_5_tmp;
reg [7:0] r25_6_tmp;
reg [7:0] r25_7_tmp;
reg [7:0] r25_8_tmp;
reg [7:0] r25_9_tmp;
reg [7:0] r25_10_tmp;
reg [7:0] r25_11_tmp;
reg [7:0] r25_12_tmp;
reg [7:0] r25_13_tmp;
reg [7:0] r25_14_tmp;
reg [7:0] r25_15_tmp;
reg [7:0] r25_16_tmp;
reg [7:0] r25_17_tmp;
reg [7:0] r25_18_tmp;
reg [7:0] r25_19_tmp;
reg [7:0] r25_20_tmp;
reg [7:0] r25_21_tmp;
reg [7:0] r25_22_tmp;
reg [7:0] r25_23_tmp;
reg [7:0] r25_24_tmp;
reg [7:0] r25_25_tmp;
reg [7:0] r25_26_tmp;
reg [7:0] r25_27_tmp;
reg [7:0] r25_28_tmp;
reg [7:0] r25_29_tmp;
reg [7:0] r25_30_tmp;
reg [7:0] r25_31_tmp;
reg [7:0] r25_32_tmp;
reg [7:0] r25_34_tmp;
reg [7:0] r25_36_tmp;
reg [7:0] r25_38_tmp;
reg [7:0] r25_41_tmp;
reg [7:0] r25_43_tmp;
reg [7:0] r25_45_tmp;
reg [7:0] r25_47_tmp;
reg [7:0] r25_48_tmp;
reg [7:0] r25_49_tmp;
reg [7:0] r25_50_tmp;
reg [7:0] r25_51_tmp;
reg [7:0] r25_52_tmp;
reg [7:0] r25_53_tmp;
reg [7:0] r25_54_tmp;
reg [7:0] r25_55_tmp;
reg [7:0] r25_56_tmp;
reg [7:0] r25_57_tmp;
reg [7:0] r25_58_tmp;
reg [7:0] r25_59_tmp;
reg [7:0] r25_60_tmp;
reg [7:0] r25_61_tmp;
reg [7:0] r25_62_tmp;
reg [7:0] r25_63_tmp;
reg [7:0] r25_64_tmp;
reg [7:0] r25_65_tmp;
reg [7:0] r25_66_tmp;
reg [7:0] r25_67_tmp;
reg [7:0] r25_68_tmp;
reg [7:0] r25_69_tmp;
reg [7:0] r25_70_tmp;
reg [7:0] r25_71_tmp;
reg [7:0] r25_72_tmp;
reg [7:0] r25_73_tmp;
reg [7:0] r25_74_tmp;
reg [7:0] r25_75_tmp;
reg [7:0] r25_76_tmp;
reg [7:0] r25_77_tmp;
reg [7:0] r25_78_tmp;
reg [7:0] r25_79_tmp;
reg [7:0] r25_80_tmp;
reg [7:0] r26_0_tmp;
reg [7:0] r26_1_tmp;
reg [7:0] r26_2_tmp;
reg [7:0] r26_3_tmp;
reg [7:0] r26_4_tmp;
reg [7:0] r26_5_tmp;
reg [7:0] r26_6_tmp;
reg [7:0] r26_7_tmp;
reg [7:0] r26_8_tmp;
reg [7:0] r26_9_tmp;
reg [7:0] r26_10_tmp;
reg [7:0] r26_11_tmp;
reg [7:0] r26_12_tmp;
reg [7:0] r26_13_tmp;
reg [7:0] r26_14_tmp;
reg [7:0] r26_15_tmp;
reg [7:0] r26_16_tmp;
reg [7:0] r26_17_tmp;
reg [7:0] r26_18_tmp;
reg [7:0] r26_19_tmp;
reg [7:0] r26_20_tmp;
reg [7:0] r26_21_tmp;
reg [7:0] r26_22_tmp;
reg [7:0] r26_23_tmp;
reg [7:0] r26_24_tmp;
reg [7:0] r26_25_tmp;
reg [7:0] r26_26_tmp;
reg [7:0] r26_27_tmp;
reg [7:0] r26_28_tmp;
reg [7:0] r26_29_tmp;
reg [7:0] r26_30_tmp;
reg [7:0] r26_31_tmp;
reg [7:0] r26_32_tmp;
reg [7:0] r26_33_tmp;
reg [7:0] r26_34_tmp;
reg [7:0] r26_35_tmp;
reg [7:0] r26_36_tmp;
reg [7:0] r26_38_tmp;
reg [7:0] r26_41_tmp;
reg [7:0] r26_43_tmp;
reg [7:0] r26_44_tmp;
reg [7:0] r26_45_tmp;
reg [7:0] r26_46_tmp;
reg [7:0] r26_47_tmp;
reg [7:0] r26_48_tmp;
reg [7:0] r26_49_tmp;
reg [7:0] r26_50_tmp;
reg [7:0] r26_51_tmp;
reg [7:0] r26_52_tmp;
reg [7:0] r26_53_tmp;
reg [7:0] r26_54_tmp;
reg [7:0] r26_55_tmp;
reg [7:0] r26_56_tmp;
reg [7:0] r26_57_tmp;
reg [7:0] r26_58_tmp;
reg [7:0] r26_59_tmp;
reg [7:0] r26_60_tmp;
reg [7:0] r26_61_tmp;
reg [7:0] r26_62_tmp;
reg [7:0] r26_63_tmp;
reg [7:0] r26_64_tmp;
reg [7:0] r26_65_tmp;
reg [7:0] r26_66_tmp;
reg [7:0] r26_67_tmp;
reg [7:0] r26_68_tmp;
reg [7:0] r26_69_tmp;
reg [7:0] r26_70_tmp;
reg [7:0] r26_71_tmp;
reg [7:0] r26_72_tmp;
reg [7:0] r26_73_tmp;
reg [7:0] r26_74_tmp;
reg [7:0] r26_75_tmp;
reg [7:0] r26_76_tmp;
reg [7:0] r26_77_tmp;
reg [7:0] r26_78_tmp;
reg [7:0] r26_79_tmp;
reg [7:0] r26_80_tmp;
reg [7:0] r27_0_tmp;
reg [7:0] r27_1_tmp;
reg [7:0] r27_2_tmp;
reg [7:0] r27_3_tmp;
reg [7:0] r27_4_tmp;
reg [7:0] r27_5_tmp;
reg [7:0] r27_6_tmp;
reg [7:0] r27_7_tmp;
reg [7:0] r27_8_tmp;
reg [7:0] r27_9_tmp;
reg [7:0] r27_10_tmp;
reg [7:0] r27_11_tmp;
reg [7:0] r27_12_tmp;
reg [7:0] r27_13_tmp;
reg [7:0] r27_14_tmp;
reg [7:0] r27_15_tmp;
reg [7:0] r27_16_tmp;
reg [7:0] r27_17_tmp;
reg [7:0] r27_18_tmp;
reg [7:0] r27_19_tmp;
reg [7:0] r27_20_tmp;
reg [7:0] r27_21_tmp;
reg [7:0] r27_22_tmp;
reg [7:0] r27_23_tmp;
reg [7:0] r27_24_tmp;
reg [7:0] r27_25_tmp;
reg [7:0] r27_26_tmp;
reg [7:0] r27_27_tmp;
reg [7:0] r27_28_tmp;
reg [7:0] r27_29_tmp;
reg [7:0] r27_30_tmp;
reg [7:0] r27_31_tmp;
reg [7:0] r27_32_tmp;
reg [7:0] r27_33_tmp;
reg [7:0] r27_34_tmp;
reg [7:0] r27_35_tmp;
reg [7:0] r27_36_tmp;
reg [7:0] r27_37_tmp;
reg [7:0] r27_38_tmp;
reg [7:0] r27_41_tmp;
reg [7:0] r27_42_tmp;
reg [7:0] r27_43_tmp;
reg [7:0] r27_44_tmp;
reg [7:0] r27_45_tmp;
reg [7:0] r27_46_tmp;
reg [7:0] r27_47_tmp;
reg [7:0] r27_48_tmp;
reg [7:0] r27_49_tmp;
reg [7:0] r27_50_tmp;
reg [7:0] r27_51_tmp;
reg [7:0] r27_52_tmp;
reg [7:0] r27_53_tmp;
reg [7:0] r27_54_tmp;
reg [7:0] r27_55_tmp;
reg [7:0] r27_56_tmp;
reg [7:0] r27_57_tmp;
reg [7:0] r27_58_tmp;
reg [7:0] r27_59_tmp;
reg [7:0] r27_60_tmp;
reg [7:0] r27_61_tmp;
reg [7:0] r27_62_tmp;
reg [7:0] r27_63_tmp;
reg [7:0] r27_64_tmp;
reg [7:0] r27_65_tmp;
reg [7:0] r27_66_tmp;
reg [7:0] r27_67_tmp;
reg [7:0] r27_68_tmp;
reg [7:0] r27_69_tmp;
reg [7:0] r27_70_tmp;
reg [7:0] r27_71_tmp;
reg [7:0] r27_72_tmp;
reg [7:0] r27_73_tmp;
reg [7:0] r27_74_tmp;
reg [7:0] r27_75_tmp;
reg [7:0] r27_76_tmp;
reg [7:0] r27_77_tmp;
reg [7:0] r27_78_tmp;
reg [7:0] r27_79_tmp;
reg [7:0] r27_80_tmp;
//-----------------------------

always @(posedge clk)begin
//--------INPUT LAYER-------------
cmp0_in0 <= x_0;
cmp0_in1 <= x_64;
r0[0] <= cmp0_out0;
r0[64] <= cmp0_out1;

cmp1_in0 <= x_1;
cmp1_in1 <= x_65;
r0[1] <= cmp1_out0;
r0[65] <= cmp1_out1;

cmp2_in0 <= x_2;
cmp2_in1 <= x_66;
r0[2] <= cmp2_out0;
r0[66] <= cmp2_out1;

cmp3_in0 <= x_3;
cmp3_in1 <= x_67;
r0[3] <= cmp3_out0;
r0[67] <= cmp3_out1;

cmp4_in0 <= x_4;
cmp4_in1 <= x_68;
r0[4] <= cmp4_out0;
r0[68] <= cmp4_out1;

cmp5_in0 <= x_5;
cmp5_in1 <= x_69;
r0[5] <= cmp5_out0;
r0[69] <= cmp5_out1;

cmp6_in0 <= x_6;
cmp6_in1 <= x_70;
r0[6] <= cmp6_out0;
r0[70] <= cmp6_out1;

cmp7_in0 <= x_7;
cmp7_in1 <= x_71;
r0[7] <= cmp7_out0;
r0[71] <= cmp7_out1;

cmp8_in0 <= x_8;
cmp8_in1 <= x_72;
r0[8] <= cmp8_out0;
r0[72] <= cmp8_out1;

cmp9_in0 <= x_9;
cmp9_in1 <= x_73;
r0[9] <= cmp9_out0;
r0[73] <= cmp9_out1;

cmp10_in0 <= x_10;
cmp10_in1 <= x_74;
r0[10] <= cmp10_out0;
r0[74] <= cmp10_out1;

cmp11_in0 <= x_11;
cmp11_in1 <= x_75;
r0[11] <= cmp11_out0;
r0[75] <= cmp11_out1;

cmp12_in0 <= x_12;
cmp12_in1 <= x_76;
r0[12] <= cmp12_out0;
r0[76] <= cmp12_out1;

cmp13_in0 <= x_13;
cmp13_in1 <= x_77;
r0[13] <= cmp13_out0;
r0[77] <= cmp13_out1;

cmp14_in0 <= x_14;
cmp14_in1 <= x_78;
r0[14] <= cmp14_out0;
r0[78] <= cmp14_out1;

cmp15_in0 <= x_15;
cmp15_in1 <= x_79;
r0[15] <= cmp15_out0;
r0[79] <= cmp15_out1;

cmp16_in0 <= x_16;
cmp16_in1 <= x_80;
r0[16] <= cmp16_out0;
r0[80] <= cmp16_out1;

r0_17_tmp <= x_17;
r0[17] <= r0_17_tmp ;
r0_18_tmp <= x_18;
r0[18] <= r0_18_tmp ;
r0_19_tmp <= x_19;
r0[19] <= r0_19_tmp ;
r0_20_tmp <= x_20;
r0[20] <= r0_20_tmp ;
r0_21_tmp <= x_21;
r0[21] <= r0_21_tmp ;
r0_22_tmp <= x_22;
r0[22] <= r0_22_tmp ;
r0_23_tmp <= x_23;
r0[23] <= r0_23_tmp ;
r0_24_tmp <= x_24;
r0[24] <= r0_24_tmp ;
r0_25_tmp <= x_25;
r0[25] <= r0_25_tmp ;
r0_26_tmp <= x_26;
r0[26] <= r0_26_tmp ;
r0_27_tmp <= x_27;
r0[27] <= r0_27_tmp ;
r0_28_tmp <= x_28;
r0[28] <= r0_28_tmp ;
r0_29_tmp <= x_29;
r0[29] <= r0_29_tmp ;
r0_30_tmp <= x_30;
r0[30] <= r0_30_tmp ;
r0_31_tmp <= x_31;
r0[31] <= r0_31_tmp ;
r0_32_tmp <= x_32;
r0[32] <= r0_32_tmp ;
r0_33_tmp <= x_33;
r0[33] <= r0_33_tmp ;
r0_34_tmp <= x_34;
r0[34] <= r0_34_tmp ;
r0_35_tmp <= x_35;
r0[35] <= r0_35_tmp ;
r0_36_tmp <= x_36;
r0[36] <= r0_36_tmp ;
r0_37_tmp <= x_37;
r0[37] <= r0_37_tmp ;
r0_38_tmp <= x_38;
r0[38] <= r0_38_tmp ;
r0_39_tmp <= x_39;
r0[39] <= r0_39_tmp ;
r0_40_tmp <= x_40;
r0[40] <= r0_40_tmp ;
r0_41_tmp <= x_41;
r0[41] <= r0_41_tmp ;
r0_42_tmp <= x_42;
r0[42] <= r0_42_tmp ;
r0_43_tmp <= x_43;
r0[43] <= r0_43_tmp ;
r0_44_tmp <= x_44;
r0[44] <= r0_44_tmp ;
r0_45_tmp <= x_45;
r0[45] <= r0_45_tmp ;
r0_46_tmp <= x_46;
r0[46] <= r0_46_tmp ;
r0_47_tmp <= x_47;
r0[47] <= r0_47_tmp ;
r0_48_tmp <= x_48;
r0[48] <= r0_48_tmp ;
r0_49_tmp <= x_49;
r0[49] <= r0_49_tmp ;
r0_50_tmp <= x_50;
r0[50] <= r0_50_tmp ;
r0_51_tmp <= x_51;
r0[51] <= r0_51_tmp ;
r0_52_tmp <= x_52;
r0[52] <= r0_52_tmp ;
r0_53_tmp <= x_53;
r0[53] <= r0_53_tmp ;
r0_54_tmp <= x_54;
r0[54] <= r0_54_tmp ;
r0_55_tmp <= x_55;
r0[55] <= r0_55_tmp ;
r0_56_tmp <= x_56;
r0[56] <= r0_56_tmp ;
r0_57_tmp <= x_57;
r0[57] <= r0_57_tmp ;
r0_58_tmp <= x_58;
r0[58] <= r0_58_tmp ;
r0_59_tmp <= x_59;
r0[59] <= r0_59_tmp ;
r0_60_tmp <= x_60;
r0[60] <= r0_60_tmp ;
r0_61_tmp <= x_61;
r0[61] <= r0_61_tmp ;
r0_62_tmp <= x_62;
r0[62] <= r0_62_tmp ;
r0_63_tmp <= x_63;
r0[63] <= r0_63_tmp ;
//--------------------------

//---------layer : 1------------
cmp17_in0 <= r0[0];
cmp17_in1 <= r0[32];
r1[0] <= cmp17_out0;
r1[32] <= cmp17_out1;

cmp18_in0 <= r0[1];
cmp18_in1 <= r0[33];
r1[1] <= cmp18_out0;
r1[33] <= cmp18_out1;

cmp19_in0 <= r0[2];
cmp19_in1 <= r0[34];
r1[2] <= cmp19_out0;
r1[34] <= cmp19_out1;

cmp20_in0 <= r0[3];
cmp20_in1 <= r0[35];
r1[3] <= cmp20_out0;
r1[35] <= cmp20_out1;

cmp21_in0 <= r0[4];
cmp21_in1 <= r0[36];
r1[4] <= cmp21_out0;
r1[36] <= cmp21_out1;

cmp22_in0 <= r0[5];
cmp22_in1 <= r0[37];
r1[5] <= cmp22_out0;
r1[37] <= cmp22_out1;

cmp23_in0 <= r0[6];
cmp23_in1 <= r0[38];
r1[6] <= cmp23_out0;
r1[38] <= cmp23_out1;

cmp24_in0 <= r0[7];
cmp24_in1 <= r0[39];
r1[7] <= cmp24_out0;
r1[39] <= cmp24_out1;

cmp25_in0 <= r0[8];
cmp25_in1 <= r0[40];
r1[8] <= cmp25_out0;
r1[40] <= cmp25_out1;

cmp26_in0 <= r0[9];
cmp26_in1 <= r0[41];
r1[9] <= cmp26_out0;
r1[41] <= cmp26_out1;

cmp27_in0 <= r0[10];
cmp27_in1 <= r0[42];
r1[10] <= cmp27_out0;
r1[42] <= cmp27_out1;

cmp28_in0 <= r0[11];
cmp28_in1 <= r0[43];
r1[11] <= cmp28_out0;
r1[43] <= cmp28_out1;

cmp29_in0 <= r0[12];
cmp29_in1 <= r0[44];
r1[12] <= cmp29_out0;
r1[44] <= cmp29_out1;

cmp30_in0 <= r0[13];
cmp30_in1 <= r0[45];
r1[13] <= cmp30_out0;
r1[45] <= cmp30_out1;

cmp31_in0 <= r0[14];
cmp31_in1 <= r0[46];
r1[14] <= cmp31_out0;
r1[46] <= cmp31_out1;

cmp32_in0 <= r0[15];
cmp32_in1 <= r0[47];
r1[15] <= cmp32_out0;
r1[47] <= cmp32_out1;

cmp33_in0 <= r0[16];
cmp33_in1 <= r0[48];
r1[16] <= cmp33_out0;
r1[48] <= cmp33_out1;

cmp34_in0 <= r0[17];
cmp34_in1 <= r0[49];
r1[17] <= cmp34_out0;
r1[49] <= cmp34_out1;

cmp35_in0 <= r0[18];
cmp35_in1 <= r0[50];
r1[18] <= cmp35_out0;
r1[50] <= cmp35_out1;

cmp36_in0 <= r0[19];
cmp36_in1 <= r0[51];
r1[19] <= cmp36_out0;
r1[51] <= cmp36_out1;

cmp37_in0 <= r0[20];
cmp37_in1 <= r0[52];
r1[20] <= cmp37_out0;
r1[52] <= cmp37_out1;

cmp38_in0 <= r0[21];
cmp38_in1 <= r0[53];
r1[21] <= cmp38_out0;
r1[53] <= cmp38_out1;

cmp39_in0 <= r0[22];
cmp39_in1 <= r0[54];
r1[22] <= cmp39_out0;
r1[54] <= cmp39_out1;

cmp40_in0 <= r0[23];
cmp40_in1 <= r0[55];
r1[23] <= cmp40_out0;
r1[55] <= cmp40_out1;

cmp41_in0 <= r0[24];
cmp41_in1 <= r0[56];
r1[24] <= cmp41_out0;
r1[56] <= cmp41_out1;

cmp42_in0 <= r0[25];
cmp42_in1 <= r0[57];
r1[25] <= cmp42_out0;
r1[57] <= cmp42_out1;

cmp43_in0 <= r0[26];
cmp43_in1 <= r0[58];
r1[26] <= cmp43_out0;
r1[58] <= cmp43_out1;

cmp44_in0 <= r0[27];
cmp44_in1 <= r0[59];
r1[27] <= cmp44_out0;
r1[59] <= cmp44_out1;

cmp45_in0 <= r0[28];
cmp45_in1 <= r0[60];
r1[28] <= cmp45_out0;
r1[60] <= cmp45_out1;

cmp46_in0 <= r0[29];
cmp46_in1 <= r0[61];
r1[29] <= cmp46_out0;
r1[61] <= cmp46_out1;

cmp47_in0 <= r0[30];
cmp47_in1 <= r0[62];
r1[30] <= cmp47_out0;
r1[62] <= cmp47_out1;

cmp48_in0 <= r0[31];
cmp48_in1 <= r0[63];
r1[31] <= cmp48_out0;
r1[63] <= cmp48_out1;

r1_64_tmp <= r0[64];
r1[64] <= r1_64_tmp;

r1_65_tmp <= r0[65];
r1[65] <= r1_65_tmp;

r1_66_tmp <= r0[66];
r1[66] <= r1_66_tmp;

r1_67_tmp <= r0[67];
r1[67] <= r1_67_tmp;

r1_68_tmp <= r0[68];
r1[68] <= r1_68_tmp;

r1_69_tmp <= r0[69];
r1[69] <= r1_69_tmp;

r1_70_tmp <= r0[70];
r1[70] <= r1_70_tmp;

r1_71_tmp <= r0[71];
r1[71] <= r1_71_tmp;

r1_72_tmp <= r0[72];
r1[72] <= r1_72_tmp;

r1_73_tmp <= r0[73];
r1[73] <= r1_73_tmp;

r1_74_tmp <= r0[74];
r1[74] <= r1_74_tmp;

r1_75_tmp <= r0[75];
r1[75] <= r1_75_tmp;

r1_76_tmp <= r0[76];
r1[76] <= r1_76_tmp;

r1_77_tmp <= r0[77];
r1[77] <= r1_77_tmp;

r1_78_tmp <= r0[78];
r1[78] <= r1_78_tmp;

r1_79_tmp <= r0[79];
r1[79] <= r1_79_tmp;

r1_80_tmp <= r0[80];
r1[80] <= r1_80_tmp;

//--------------------------
//---------layer : 2------------
cmp49_in0 <= r1[32];
cmp49_in1 <= r1[64];
r2[32] <= cmp49_out0;
r2[64] <= cmp49_out1;

cmp50_in0 <= r1[33];
cmp50_in1 <= r1[65];
r2[33] <= cmp50_out0;
r2[65] <= cmp50_out1;

cmp51_in0 <= r1[34];
cmp51_in1 <= r1[66];
r2[34] <= cmp51_out0;
r2[66] <= cmp51_out1;

cmp52_in0 <= r1[35];
cmp52_in1 <= r1[67];
r2[35] <= cmp52_out0;
r2[67] <= cmp52_out1;

cmp53_in0 <= r1[36];
cmp53_in1 <= r1[68];
r2[36] <= cmp53_out0;
r2[68] <= cmp53_out1;

cmp54_in0 <= r1[37];
cmp54_in1 <= r1[69];
r2[37] <= cmp54_out0;
r2[69] <= cmp54_out1;

cmp55_in0 <= r1[38];
cmp55_in1 <= r1[70];
r2[38] <= cmp55_out0;
r2[70] <= cmp55_out1;

cmp56_in0 <= r1[39];
cmp56_in1 <= r1[71];
r2[39] <= cmp56_out0;
r2[71] <= cmp56_out1;

cmp57_in0 <= r1[40];
cmp57_in1 <= r1[72];
r2[40] <= cmp57_out0;
r2[72] <= cmp57_out1;

cmp58_in0 <= r1[41];
cmp58_in1 <= r1[73];
r2[41] <= cmp58_out0;
r2[73] <= cmp58_out1;

cmp59_in0 <= r1[42];
cmp59_in1 <= r1[74];
r2[42] <= cmp59_out0;
r2[74] <= cmp59_out1;

cmp60_in0 <= r1[43];
cmp60_in1 <= r1[75];
r2[43] <= cmp60_out0;
r2[75] <= cmp60_out1;

cmp61_in0 <= r1[44];
cmp61_in1 <= r1[76];
r2[44] <= cmp61_out0;
r2[76] <= cmp61_out1;

cmp62_in0 <= r1[45];
cmp62_in1 <= r1[77];
r2[45] <= cmp62_out0;
r2[77] <= cmp62_out1;

cmp63_in0 <= r1[46];
cmp63_in1 <= r1[78];
r2[46] <= cmp63_out0;
r2[78] <= cmp63_out1;

cmp64_in0 <= r1[47];
cmp64_in1 <= r1[79];
r2[47] <= cmp64_out0;
r2[79] <= cmp64_out1;

cmp65_in0 <= r1[48];
cmp65_in1 <= r1[80];
r2[48] <= cmp65_out0;
r2[80] <= cmp65_out1;

cmp66_in0 <= r1[0];
cmp66_in1 <= r1[16];
r2[0] <= cmp66_out0;
r2[16] <= cmp66_out1;

cmp67_in0 <= r1[1];
cmp67_in1 <= r1[17];
r2[1] <= cmp67_out0;
r2[17] <= cmp67_out1;

cmp68_in0 <= r1[2];
cmp68_in1 <= r1[18];
r2[2] <= cmp68_out0;
r2[18] <= cmp68_out1;

cmp69_in0 <= r1[3];
cmp69_in1 <= r1[19];
r2[3] <= cmp69_out0;
r2[19] <= cmp69_out1;

cmp70_in0 <= r1[4];
cmp70_in1 <= r1[20];
r2[4] <= cmp70_out0;
r2[20] <= cmp70_out1;

cmp71_in0 <= r1[5];
cmp71_in1 <= r1[21];
r2[5] <= cmp71_out0;
r2[21] <= cmp71_out1;

cmp72_in0 <= r1[6];
cmp72_in1 <= r1[22];
r2[6] <= cmp72_out0;
r2[22] <= cmp72_out1;

cmp73_in0 <= r1[7];
cmp73_in1 <= r1[23];
r2[7] <= cmp73_out0;
r2[23] <= cmp73_out1;

cmp74_in0 <= r1[8];
cmp74_in1 <= r1[24];
r2[8] <= cmp74_out0;
r2[24] <= cmp74_out1;

cmp75_in0 <= r1[9];
cmp75_in1 <= r1[25];
r2[9] <= cmp75_out0;
r2[25] <= cmp75_out1;

cmp76_in0 <= r1[10];
cmp76_in1 <= r1[26];
r2[10] <= cmp76_out0;
r2[26] <= cmp76_out1;

cmp77_in0 <= r1[11];
cmp77_in1 <= r1[27];
r2[11] <= cmp77_out0;
r2[27] <= cmp77_out1;

cmp78_in0 <= r1[12];
cmp78_in1 <= r1[28];
r2[12] <= cmp78_out0;
r2[28] <= cmp78_out1;

cmp79_in0 <= r1[13];
cmp79_in1 <= r1[29];
r2[13] <= cmp79_out0;
r2[29] <= cmp79_out1;

cmp80_in0 <= r1[14];
cmp80_in1 <= r1[30];
r2[14] <= cmp80_out0;
r2[30] <= cmp80_out1;

cmp81_in0 <= r1[15];
cmp81_in1 <= r1[31];
r2[15] <= cmp81_out0;
r2[31] <= cmp81_out1;

r2_49_tmp <= r1[49];
r2[49] <= r2_49_tmp;

r2_50_tmp <= r1[50];
r2[50] <= r2_50_tmp;

r2_51_tmp <= r1[51];
r2[51] <= r2_51_tmp;

r2_52_tmp <= r1[52];
r2[52] <= r2_52_tmp;

r2_53_tmp <= r1[53];
r2[53] <= r2_53_tmp;

r2_54_tmp <= r1[54];
r2[54] <= r2_54_tmp;

r2_55_tmp <= r1[55];
r2[55] <= r2_55_tmp;

r2_56_tmp <= r1[56];
r2[56] <= r2_56_tmp;

r2_57_tmp <= r1[57];
r2[57] <= r2_57_tmp;

r2_58_tmp <= r1[58];
r2[58] <= r2_58_tmp;

r2_59_tmp <= r1[59];
r2[59] <= r2_59_tmp;

r2_60_tmp <= r1[60];
r2[60] <= r2_60_tmp;

r2_61_tmp <= r1[61];
r2[61] <= r2_61_tmp;

r2_62_tmp <= r1[62];
r2[62] <= r2_62_tmp;

r2_63_tmp <= r1[63];
r2[63] <= r2_63_tmp;

//--------------------------
//---------layer : 3------------
cmp82_in0 <= r2[32];
cmp82_in1 <= r2[48];
r3[32] <= cmp82_out0;
r3[48] <= cmp82_out1;

cmp83_in0 <= r2[33];
cmp83_in1 <= r2[49];
r3[33] <= cmp83_out0;
r3[49] <= cmp83_out1;

cmp84_in0 <= r2[34];
cmp84_in1 <= r2[50];
r3[34] <= cmp84_out0;
r3[50] <= cmp84_out1;

cmp85_in0 <= r2[35];
cmp85_in1 <= r2[51];
r3[35] <= cmp85_out0;
r3[51] <= cmp85_out1;

cmp86_in0 <= r2[36];
cmp86_in1 <= r2[52];
r3[36] <= cmp86_out0;
r3[52] <= cmp86_out1;

cmp87_in0 <= r2[37];
cmp87_in1 <= r2[53];
r3[37] <= cmp87_out0;
r3[53] <= cmp87_out1;

cmp88_in0 <= r2[38];
cmp88_in1 <= r2[54];
r3[38] <= cmp88_out0;
r3[54] <= cmp88_out1;

cmp89_in0 <= r2[39];
cmp89_in1 <= r2[55];
r3[39] <= cmp89_out0;
r3[55] <= cmp89_out1;

cmp90_in0 <= r2[40];
cmp90_in1 <= r2[56];
r3[40] <= cmp90_out0;
r3[56] <= cmp90_out1;

cmp91_in0 <= r2[41];
cmp91_in1 <= r2[57];
r3[41] <= cmp91_out0;
r3[57] <= cmp91_out1;

cmp92_in0 <= r2[42];
cmp92_in1 <= r2[58];
r3[42] <= cmp92_out0;
r3[58] <= cmp92_out1;

cmp93_in0 <= r2[43];
cmp93_in1 <= r2[59];
r3[43] <= cmp93_out0;
r3[59] <= cmp93_out1;

cmp94_in0 <= r2[44];
cmp94_in1 <= r2[60];
r3[44] <= cmp94_out0;
r3[60] <= cmp94_out1;

cmp95_in0 <= r2[45];
cmp95_in1 <= r2[61];
r3[45] <= cmp95_out0;
r3[61] <= cmp95_out1;

cmp96_in0 <= r2[46];
cmp96_in1 <= r2[62];
r3[46] <= cmp96_out0;
r3[62] <= cmp96_out1;

cmp97_in0 <= r2[47];
cmp97_in1 <= r2[63];
r3[47] <= cmp97_out0;
r3[63] <= cmp97_out1;

cmp98_in0 <= r2[64];
cmp98_in1 <= r2[80];
r3[64] <= cmp98_out0;
r3[80] <= cmp98_out1;

r3_0_tmp <= r2[0];
r3[0] <= r3_0_tmp;

r3_1_tmp <= r2[1];
r3[1] <= r3_1_tmp;

r3_2_tmp <= r2[2];
r3[2] <= r3_2_tmp;

r3_3_tmp <= r2[3];
r3[3] <= r3_3_tmp;

r3_4_tmp <= r2[4];
r3[4] <= r3_4_tmp;

r3_5_tmp <= r2[5];
r3[5] <= r3_5_tmp;

r3_6_tmp <= r2[6];
r3[6] <= r3_6_tmp;

r3_7_tmp <= r2[7];
r3[7] <= r3_7_tmp;

r3_8_tmp <= r2[8];
r3[8] <= r3_8_tmp;

r3_9_tmp <= r2[9];
r3[9] <= r3_9_tmp;

r3_10_tmp <= r2[10];
r3[10] <= r3_10_tmp;

r3_11_tmp <= r2[11];
r3[11] <= r3_11_tmp;

r3_12_tmp <= r2[12];
r3[12] <= r3_12_tmp;

r3_13_tmp <= r2[13];
r3[13] <= r3_13_tmp;

r3_14_tmp <= r2[14];
r3[14] <= r3_14_tmp;

r3_15_tmp <= r2[15];
r3[15] <= r3_15_tmp;

r3_16_tmp <= r2[16];
r3[16] <= r3_16_tmp;

r3_17_tmp <= r2[17];
r3[17] <= r3_17_tmp;

r3_18_tmp <= r2[18];
r3[18] <= r3_18_tmp;

r3_19_tmp <= r2[19];
r3[19] <= r3_19_tmp;

r3_20_tmp <= r2[20];
r3[20] <= r3_20_tmp;

r3_21_tmp <= r2[21];
r3[21] <= r3_21_tmp;

r3_22_tmp <= r2[22];
r3[22] <= r3_22_tmp;

r3_23_tmp <= r2[23];
r3[23] <= r3_23_tmp;

r3_24_tmp <= r2[24];
r3[24] <= r3_24_tmp;

r3_25_tmp <= r2[25];
r3[25] <= r3_25_tmp;

r3_26_tmp <= r2[26];
r3[26] <= r3_26_tmp;

r3_27_tmp <= r2[27];
r3[27] <= r3_27_tmp;

r3_28_tmp <= r2[28];
r3[28] <= r3_28_tmp;

r3_29_tmp <= r2[29];
r3[29] <= r3_29_tmp;

r3_30_tmp <= r2[30];
r3[30] <= r3_30_tmp;

r3_31_tmp <= r2[31];
r3[31] <= r3_31_tmp;

r3_65_tmp <= r2[65];
r3[65] <= r3_65_tmp;

r3_66_tmp <= r2[66];
r3[66] <= r3_66_tmp;

r3_67_tmp <= r2[67];
r3[67] <= r3_67_tmp;

r3_68_tmp <= r2[68];
r3[68] <= r3_68_tmp;

r3_69_tmp <= r2[69];
r3[69] <= r3_69_tmp;

r3_70_tmp <= r2[70];
r3[70] <= r3_70_tmp;

r3_71_tmp <= r2[71];
r3[71] <= r3_71_tmp;

r3_72_tmp <= r2[72];
r3[72] <= r3_72_tmp;

r3_73_tmp <= r2[73];
r3[73] <= r3_73_tmp;

r3_74_tmp <= r2[74];
r3[74] <= r3_74_tmp;

r3_75_tmp <= r2[75];
r3[75] <= r3_75_tmp;

r3_76_tmp <= r2[76];
r3[76] <= r3_76_tmp;

r3_77_tmp <= r2[77];
r3[77] <= r3_77_tmp;

r3_78_tmp <= r2[78];
r3[78] <= r3_78_tmp;

r3_79_tmp <= r2[79];
r3[79] <= r3_79_tmp;

//--------------------------
//---------layer : 4------------
cmp99_in0 <= r3[16];
cmp99_in1 <= r3[64];
r4[16] <= cmp99_out0;
r4[64] <= cmp99_out1;

cmp100_in0 <= r3[17];
cmp100_in1 <= r3[65];
r4[17] <= cmp100_out0;
r4[65] <= cmp100_out1;

cmp101_in0 <= r3[18];
cmp101_in1 <= r3[66];
r4[18] <= cmp101_out0;
r4[66] <= cmp101_out1;

cmp102_in0 <= r3[19];
cmp102_in1 <= r3[67];
r4[19] <= cmp102_out0;
r4[67] <= cmp102_out1;

cmp103_in0 <= r3[20];
cmp103_in1 <= r3[68];
r4[20] <= cmp103_out0;
r4[68] <= cmp103_out1;

cmp104_in0 <= r3[21];
cmp104_in1 <= r3[69];
r4[21] <= cmp104_out0;
r4[69] <= cmp104_out1;

cmp105_in0 <= r3[22];
cmp105_in1 <= r3[70];
r4[22] <= cmp105_out0;
r4[70] <= cmp105_out1;

cmp106_in0 <= r3[23];
cmp106_in1 <= r3[71];
r4[23] <= cmp106_out0;
r4[71] <= cmp106_out1;

cmp107_in0 <= r3[24];
cmp107_in1 <= r3[72];
r4[24] <= cmp107_out0;
r4[72] <= cmp107_out1;

cmp108_in0 <= r3[25];
cmp108_in1 <= r3[73];
r4[25] <= cmp108_out0;
r4[73] <= cmp108_out1;

cmp109_in0 <= r3[26];
cmp109_in1 <= r3[74];
r4[26] <= cmp109_out0;
r4[74] <= cmp109_out1;

cmp110_in0 <= r3[27];
cmp110_in1 <= r3[75];
r4[27] <= cmp110_out0;
r4[75] <= cmp110_out1;

cmp111_in0 <= r3[28];
cmp111_in1 <= r3[76];
r4[28] <= cmp111_out0;
r4[76] <= cmp111_out1;

cmp112_in0 <= r3[29];
cmp112_in1 <= r3[77];
r4[29] <= cmp112_out0;
r4[77] <= cmp112_out1;

cmp113_in0 <= r3[30];
cmp113_in1 <= r3[78];
r4[30] <= cmp113_out0;
r4[78] <= cmp113_out1;

cmp114_in0 <= r3[31];
cmp114_in1 <= r3[79];
r4[31] <= cmp114_out0;
r4[79] <= cmp114_out1;

r4_0_tmp <= r3[0];
r4[0] <= r4_0_tmp;

r4_1_tmp <= r3[1];
r4[1] <= r4_1_tmp;

r4_2_tmp <= r3[2];
r4[2] <= r4_2_tmp;

r4_3_tmp <= r3[3];
r4[3] <= r4_3_tmp;

r4_4_tmp <= r3[4];
r4[4] <= r4_4_tmp;

r4_5_tmp <= r3[5];
r4[5] <= r4_5_tmp;

r4_6_tmp <= r3[6];
r4[6] <= r4_6_tmp;

r4_7_tmp <= r3[7];
r4[7] <= r4_7_tmp;

r4_8_tmp <= r3[8];
r4[8] <= r4_8_tmp;

r4_9_tmp <= r3[9];
r4[9] <= r4_9_tmp;

r4_10_tmp <= r3[10];
r4[10] <= r4_10_tmp;

r4_11_tmp <= r3[11];
r4[11] <= r4_11_tmp;

r4_12_tmp <= r3[12];
r4[12] <= r4_12_tmp;

r4_13_tmp <= r3[13];
r4[13] <= r4_13_tmp;

r4_14_tmp <= r3[14];
r4[14] <= r4_14_tmp;

r4_15_tmp <= r3[15];
r4[15] <= r4_15_tmp;

r4_32_tmp <= r3[32];
r4[32] <= r4_32_tmp;

r4_33_tmp <= r3[33];
r4[33] <= r4_33_tmp;

r4_34_tmp <= r3[34];
r4[34] <= r4_34_tmp;

r4_35_tmp <= r3[35];
r4[35] <= r4_35_tmp;

r4_36_tmp <= r3[36];
r4[36] <= r4_36_tmp;

r4_37_tmp <= r3[37];
r4[37] <= r4_37_tmp;

r4_38_tmp <= r3[38];
r4[38] <= r4_38_tmp;

r4_39_tmp <= r3[39];
r4[39] <= r4_39_tmp;

r4_40_tmp <= r3[40];
r4[40] <= r4_40_tmp;

r4_41_tmp <= r3[41];
r4[41] <= r4_41_tmp;

r4_42_tmp <= r3[42];
r4[42] <= r4_42_tmp;

r4_43_tmp <= r3[43];
r4[43] <= r4_43_tmp;

r4_44_tmp <= r3[44];
r4[44] <= r4_44_tmp;

r4_45_tmp <= r3[45];
r4[45] <= r4_45_tmp;

r4_46_tmp <= r3[46];
r4[46] <= r4_46_tmp;

r4_47_tmp <= r3[47];
r4[47] <= r4_47_tmp;

r4_48_tmp <= r3[48];
r4[48] <= r4_48_tmp;

r4_49_tmp <= r3[49];
r4[49] <= r4_49_tmp;

r4_50_tmp <= r3[50];
r4[50] <= r4_50_tmp;

r4_51_tmp <= r3[51];
r4[51] <= r4_51_tmp;

r4_52_tmp <= r3[52];
r4[52] <= r4_52_tmp;

r4_53_tmp <= r3[53];
r4[53] <= r4_53_tmp;

r4_54_tmp <= r3[54];
r4[54] <= r4_54_tmp;

r4_55_tmp <= r3[55];
r4[55] <= r4_55_tmp;

r4_56_tmp <= r3[56];
r4[56] <= r4_56_tmp;

r4_57_tmp <= r3[57];
r4[57] <= r4_57_tmp;

r4_58_tmp <= r3[58];
r4[58] <= r4_58_tmp;

r4_59_tmp <= r3[59];
r4[59] <= r4_59_tmp;

r4_60_tmp <= r3[60];
r4[60] <= r4_60_tmp;

r4_61_tmp <= r3[61];
r4[61] <= r4_61_tmp;

r4_62_tmp <= r3[62];
r4[62] <= r4_62_tmp;

r4_63_tmp <= r3[63];
r4[63] <= r4_63_tmp;

r4_80_tmp <= r3[80];
r4[80] <= r4_80_tmp;

//--------------------------
//---------layer : 5------------
cmp115_in0 <= r4[16];
cmp115_in1 <= r4[32];
r5[16] <= cmp115_out0;
r5[32] <= cmp115_out1;

cmp116_in0 <= r4[17];
cmp116_in1 <= r4[33];
r5[17] <= cmp116_out0;
r5[33] <= cmp116_out1;

cmp117_in0 <= r4[18];
cmp117_in1 <= r4[34];
r5[18] <= cmp117_out0;
r5[34] <= cmp117_out1;

cmp118_in0 <= r4[19];
cmp118_in1 <= r4[35];
r5[19] <= cmp118_out0;
r5[35] <= cmp118_out1;

cmp119_in0 <= r4[20];
cmp119_in1 <= r4[36];
r5[20] <= cmp119_out0;
r5[36] <= cmp119_out1;

cmp120_in0 <= r4[21];
cmp120_in1 <= r4[37];
r5[21] <= cmp120_out0;
r5[37] <= cmp120_out1;

cmp121_in0 <= r4[22];
cmp121_in1 <= r4[38];
r5[22] <= cmp121_out0;
r5[38] <= cmp121_out1;

cmp122_in0 <= r4[23];
cmp122_in1 <= r4[39];
r5[23] <= cmp122_out0;
r5[39] <= cmp122_out1;

cmp123_in0 <= r4[24];
cmp123_in1 <= r4[40];
r5[24] <= cmp123_out0;
r5[40] <= cmp123_out1;

cmp124_in0 <= r4[25];
cmp124_in1 <= r4[41];
r5[25] <= cmp124_out0;
r5[41] <= cmp124_out1;

cmp125_in0 <= r4[26];
cmp125_in1 <= r4[42];
r5[26] <= cmp125_out0;
r5[42] <= cmp125_out1;

cmp126_in0 <= r4[27];
cmp126_in1 <= r4[43];
r5[27] <= cmp126_out0;
r5[43] <= cmp126_out1;

cmp127_in0 <= r4[28];
cmp127_in1 <= r4[44];
r5[28] <= cmp127_out0;
r5[44] <= cmp127_out1;

cmp128_in0 <= r4[29];
cmp128_in1 <= r4[45];
r5[29] <= cmp128_out0;
r5[45] <= cmp128_out1;

cmp129_in0 <= r4[30];
cmp129_in1 <= r4[46];
r5[30] <= cmp129_out0;
r5[46] <= cmp129_out1;

cmp130_in0 <= r4[31];
cmp130_in1 <= r4[47];
r5[31] <= cmp130_out0;
r5[47] <= cmp130_out1;

cmp131_in0 <= r4[48];
cmp131_in1 <= r4[64];
r5[48] <= cmp131_out0;
r5[64] <= cmp131_out1;

cmp132_in0 <= r4[49];
cmp132_in1 <= r4[65];
r5[49] <= cmp132_out0;
r5[65] <= cmp132_out1;

cmp133_in0 <= r4[50];
cmp133_in1 <= r4[66];
r5[50] <= cmp133_out0;
r5[66] <= cmp133_out1;

cmp134_in0 <= r4[51];
cmp134_in1 <= r4[67];
r5[51] <= cmp134_out0;
r5[67] <= cmp134_out1;

cmp135_in0 <= r4[52];
cmp135_in1 <= r4[68];
r5[52] <= cmp135_out0;
r5[68] <= cmp135_out1;

cmp136_in0 <= r4[53];
cmp136_in1 <= r4[69];
r5[53] <= cmp136_out0;
r5[69] <= cmp136_out1;

cmp137_in0 <= r4[54];
cmp137_in1 <= r4[70];
r5[54] <= cmp137_out0;
r5[70] <= cmp137_out1;

cmp138_in0 <= r4[55];
cmp138_in1 <= r4[71];
r5[55] <= cmp138_out0;
r5[71] <= cmp138_out1;

cmp139_in0 <= r4[56];
cmp139_in1 <= r4[72];
r5[56] <= cmp139_out0;
r5[72] <= cmp139_out1;

cmp140_in0 <= r4[57];
cmp140_in1 <= r4[73];
r5[57] <= cmp140_out0;
r5[73] <= cmp140_out1;

cmp141_in0 <= r4[58];
cmp141_in1 <= r4[74];
r5[58] <= cmp141_out0;
r5[74] <= cmp141_out1;

cmp142_in0 <= r4[59];
cmp142_in1 <= r4[75];
r5[59] <= cmp142_out0;
r5[75] <= cmp142_out1;

cmp143_in0 <= r4[60];
cmp143_in1 <= r4[76];
r5[60] <= cmp143_out0;
r5[76] <= cmp143_out1;

cmp144_in0 <= r4[61];
cmp144_in1 <= r4[77];
r5[61] <= cmp144_out0;
r5[77] <= cmp144_out1;

cmp145_in0 <= r4[62];
cmp145_in1 <= r4[78];
r5[62] <= cmp145_out0;
r5[78] <= cmp145_out1;

cmp146_in0 <= r4[63];
cmp146_in1 <= r4[79];
r5[63] <= cmp146_out0;
r5[79] <= cmp146_out1;

cmp147_in0 <= r4[0];
cmp147_in1 <= r4[8];
r5[0] <= cmp147_out0;
r5[8] <= cmp147_out1;

cmp148_in0 <= r4[1];
cmp148_in1 <= r4[9];
r5[1] <= cmp148_out0;
r5[9] <= cmp148_out1;

cmp149_in0 <= r4[2];
cmp149_in1 <= r4[10];
r5[2] <= cmp149_out0;
r5[10] <= cmp149_out1;

cmp150_in0 <= r4[3];
cmp150_in1 <= r4[11];
r5[3] <= cmp150_out0;
r5[11] <= cmp150_out1;

cmp151_in0 <= r4[4];
cmp151_in1 <= r4[12];
r5[4] <= cmp151_out0;
r5[12] <= cmp151_out1;

cmp152_in0 <= r4[5];
cmp152_in1 <= r4[13];
r5[5] <= cmp152_out0;
r5[13] <= cmp152_out1;

cmp153_in0 <= r4[6];
cmp153_in1 <= r4[14];
r5[6] <= cmp153_out0;
r5[14] <= cmp153_out1;

cmp154_in0 <= r4[7];
cmp154_in1 <= r4[15];
r5[7] <= cmp154_out0;
r5[15] <= cmp154_out1;

r5_80_tmp <= r4[80];
r5[80] <= r5_80_tmp;

//--------------------------
//---------layer : 6------------
cmp155_in0 <= r5[16];
cmp155_in1 <= r5[24];
r6[16] <= cmp155_out0;
r6[24] <= cmp155_out1;

cmp156_in0 <= r5[17];
cmp156_in1 <= r5[25];
r6[17] <= cmp156_out0;
r6[25] <= cmp156_out1;

cmp157_in0 <= r5[18];
cmp157_in1 <= r5[26];
r6[18] <= cmp157_out0;
r6[26] <= cmp157_out1;

cmp158_in0 <= r5[19];
cmp158_in1 <= r5[27];
r6[19] <= cmp158_out0;
r6[27] <= cmp158_out1;

cmp159_in0 <= r5[20];
cmp159_in1 <= r5[28];
r6[20] <= cmp159_out0;
r6[28] <= cmp159_out1;

cmp160_in0 <= r5[21];
cmp160_in1 <= r5[29];
r6[21] <= cmp160_out0;
r6[29] <= cmp160_out1;

cmp161_in0 <= r5[22];
cmp161_in1 <= r5[30];
r6[22] <= cmp161_out0;
r6[30] <= cmp161_out1;

cmp162_in0 <= r5[23];
cmp162_in1 <= r5[31];
r6[23] <= cmp162_out0;
r6[31] <= cmp162_out1;

cmp163_in0 <= r5[32];
cmp163_in1 <= r5[40];
r6[32] <= cmp163_out0;
r6[40] <= cmp163_out1;

cmp164_in0 <= r5[33];
cmp164_in1 <= r5[41];
r6[33] <= cmp164_out0;
r6[41] <= cmp164_out1;

cmp165_in0 <= r5[34];
cmp165_in1 <= r5[42];
r6[34] <= cmp165_out0;
r6[42] <= cmp165_out1;

cmp166_in0 <= r5[35];
cmp166_in1 <= r5[43];
r6[35] <= cmp166_out0;
r6[43] <= cmp166_out1;

cmp167_in0 <= r5[36];
cmp167_in1 <= r5[44];
r6[36] <= cmp167_out0;
r6[44] <= cmp167_out1;

cmp168_in0 <= r5[37];
cmp168_in1 <= r5[45];
r6[37] <= cmp168_out0;
r6[45] <= cmp168_out1;

cmp169_in0 <= r5[38];
cmp169_in1 <= r5[46];
r6[38] <= cmp169_out0;
r6[46] <= cmp169_out1;

cmp170_in0 <= r5[39];
cmp170_in1 <= r5[47];
r6[39] <= cmp170_out0;
r6[47] <= cmp170_out1;

cmp171_in0 <= r5[48];
cmp171_in1 <= r5[56];
r6[48] <= cmp171_out0;
r6[56] <= cmp171_out1;

cmp172_in0 <= r5[49];
cmp172_in1 <= r5[57];
r6[49] <= cmp172_out0;
r6[57] <= cmp172_out1;

cmp173_in0 <= r5[50];
cmp173_in1 <= r5[58];
r6[50] <= cmp173_out0;
r6[58] <= cmp173_out1;

cmp174_in0 <= r5[51];
cmp174_in1 <= r5[59];
r6[51] <= cmp174_out0;
r6[59] <= cmp174_out1;

cmp175_in0 <= r5[52];
cmp175_in1 <= r5[60];
r6[52] <= cmp175_out0;
r6[60] <= cmp175_out1;

cmp176_in0 <= r5[53];
cmp176_in1 <= r5[61];
r6[53] <= cmp176_out0;
r6[61] <= cmp176_out1;

cmp177_in0 <= r5[54];
cmp177_in1 <= r5[62];
r6[54] <= cmp177_out0;
r6[62] <= cmp177_out1;

cmp178_in0 <= r5[55];
cmp178_in1 <= r5[63];
r6[55] <= cmp178_out0;
r6[63] <= cmp178_out1;

cmp179_in0 <= r5[64];
cmp179_in1 <= r5[72];
r6[64] <= cmp179_out0;
r6[72] <= cmp179_out1;

cmp180_in0 <= r5[65];
cmp180_in1 <= r5[73];
r6[65] <= cmp180_out0;
r6[73] <= cmp180_out1;

cmp181_in0 <= r5[66];
cmp181_in1 <= r5[74];
r6[66] <= cmp181_out0;
r6[74] <= cmp181_out1;

cmp182_in0 <= r5[67];
cmp182_in1 <= r5[75];
r6[67] <= cmp182_out0;
r6[75] <= cmp182_out1;

cmp183_in0 <= r5[68];
cmp183_in1 <= r5[76];
r6[68] <= cmp183_out0;
r6[76] <= cmp183_out1;

cmp184_in0 <= r5[69];
cmp184_in1 <= r5[77];
r6[69] <= cmp184_out0;
r6[77] <= cmp184_out1;

cmp185_in0 <= r5[70];
cmp185_in1 <= r5[78];
r6[70] <= cmp185_out0;
r6[78] <= cmp185_out1;

cmp186_in0 <= r5[71];
cmp186_in1 <= r5[79];
r6[71] <= cmp186_out0;
r6[79] <= cmp186_out1;

r6_0_tmp <= r5[0];
r6[0] <= r6_0_tmp;

r6_1_tmp <= r5[1];
r6[1] <= r6_1_tmp;

r6_2_tmp <= r5[2];
r6[2] <= r6_2_tmp;

r6_3_tmp <= r5[3];
r6[3] <= r6_3_tmp;

r6_4_tmp <= r5[4];
r6[4] <= r6_4_tmp;

r6_5_tmp <= r5[5];
r6[5] <= r6_5_tmp;

r6_6_tmp <= r5[6];
r6[6] <= r6_6_tmp;

r6_7_tmp <= r5[7];
r6[7] <= r6_7_tmp;

r6_8_tmp <= r5[8];
r6[8] <= r6_8_tmp;

r6_9_tmp <= r5[9];
r6[9] <= r6_9_tmp;

r6_10_tmp <= r5[10];
r6[10] <= r6_10_tmp;

r6_11_tmp <= r5[11];
r6[11] <= r6_11_tmp;

r6_12_tmp <= r5[12];
r6[12] <= r6_12_tmp;

r6_13_tmp <= r5[13];
r6[13] <= r6_13_tmp;

r6_14_tmp <= r5[14];
r6[14] <= r6_14_tmp;

r6_15_tmp <= r5[15];
r6[15] <= r6_15_tmp;

r6_80_tmp <= r5[80];
r6[80] <= r6_80_tmp;

//--------------------------
//---------layer : 7------------
cmp187_in0 <= r6[8];
cmp187_in1 <= r6[64];
r7[8] <= cmp187_out0;
r7[64] <= cmp187_out1;

cmp188_in0 <= r6[9];
cmp188_in1 <= r6[65];
r7[9] <= cmp188_out0;
r7[65] <= cmp188_out1;

cmp189_in0 <= r6[10];
cmp189_in1 <= r6[66];
r7[10] <= cmp189_out0;
r7[66] <= cmp189_out1;

cmp190_in0 <= r6[11];
cmp190_in1 <= r6[67];
r7[11] <= cmp190_out0;
r7[67] <= cmp190_out1;

cmp191_in0 <= r6[12];
cmp191_in1 <= r6[68];
r7[12] <= cmp191_out0;
r7[68] <= cmp191_out1;

cmp192_in0 <= r6[13];
cmp192_in1 <= r6[69];
r7[13] <= cmp192_out0;
r7[69] <= cmp192_out1;

cmp193_in0 <= r6[14];
cmp193_in1 <= r6[70];
r7[14] <= cmp193_out0;
r7[70] <= cmp193_out1;

cmp194_in0 <= r6[15];
cmp194_in1 <= r6[71];
r7[15] <= cmp194_out0;
r7[71] <= cmp194_out1;

cmp195_in0 <= r6[24];
cmp195_in1 <= r6[80];
r7[24] <= cmp195_out0;
r7[80] <= cmp195_out1;

r7_0_tmp <= r6[0];
r7[0] <= r7_0_tmp;

r7_1_tmp <= r6[1];
r7[1] <= r7_1_tmp;

r7_2_tmp <= r6[2];
r7[2] <= r7_2_tmp;

r7_3_tmp <= r6[3];
r7[3] <= r7_3_tmp;

r7_4_tmp <= r6[4];
r7[4] <= r7_4_tmp;

r7_5_tmp <= r6[5];
r7[5] <= r7_5_tmp;

r7_6_tmp <= r6[6];
r7[6] <= r7_6_tmp;

r7_7_tmp <= r6[7];
r7[7] <= r7_7_tmp;

r7_16_tmp <= r6[16];
r7[16] <= r7_16_tmp;

r7_17_tmp <= r6[17];
r7[17] <= r7_17_tmp;

r7_18_tmp <= r6[18];
r7[18] <= r7_18_tmp;

r7_19_tmp <= r6[19];
r7[19] <= r7_19_tmp;

r7_20_tmp <= r6[20];
r7[20] <= r7_20_tmp;

r7_21_tmp <= r6[21];
r7[21] <= r7_21_tmp;

r7_22_tmp <= r6[22];
r7[22] <= r7_22_tmp;

r7_23_tmp <= r6[23];
r7[23] <= r7_23_tmp;

r7_25_tmp <= r6[25];
r7[25] <= r7_25_tmp;

r7_26_tmp <= r6[26];
r7[26] <= r7_26_tmp;

r7_27_tmp <= r6[27];
r7[27] <= r7_27_tmp;

r7_28_tmp <= r6[28];
r7[28] <= r7_28_tmp;

r7_29_tmp <= r6[29];
r7[29] <= r7_29_tmp;

r7_30_tmp <= r6[30];
r7[30] <= r7_30_tmp;

r7_31_tmp <= r6[31];
r7[31] <= r7_31_tmp;

r7_32_tmp <= r6[32];
r7[32] <= r7_32_tmp;

r7_33_tmp <= r6[33];
r7[33] <= r7_33_tmp;

r7_34_tmp <= r6[34];
r7[34] <= r7_34_tmp;

r7_35_tmp <= r6[35];
r7[35] <= r7_35_tmp;

r7_36_tmp <= r6[36];
r7[36] <= r7_36_tmp;

r7_37_tmp <= r6[37];
r7[37] <= r7_37_tmp;

r7_38_tmp <= r6[38];
r7[38] <= r7_38_tmp;

r7_39_tmp <= r6[39];
r7[39] <= r7_39_tmp;

r7_40_tmp <= r6[40];
r7[40] <= r7_40_tmp;

r7_41_tmp <= r6[41];
r7[41] <= r7_41_tmp;

r7_42_tmp <= r6[42];
r7[42] <= r7_42_tmp;

r7_43_tmp <= r6[43];
r7[43] <= r7_43_tmp;

r7_44_tmp <= r6[44];
r7[44] <= r7_44_tmp;

r7_45_tmp <= r6[45];
r7[45] <= r7_45_tmp;

r7_46_tmp <= r6[46];
r7[46] <= r7_46_tmp;

r7_47_tmp <= r6[47];
r7[47] <= r7_47_tmp;

r7_48_tmp <= r6[48];
r7[48] <= r7_48_tmp;

r7_49_tmp <= r6[49];
r7[49] <= r7_49_tmp;

r7_50_tmp <= r6[50];
r7[50] <= r7_50_tmp;

r7_51_tmp <= r6[51];
r7[51] <= r7_51_tmp;

r7_52_tmp <= r6[52];
r7[52] <= r7_52_tmp;

r7_53_tmp <= r6[53];
r7[53] <= r7_53_tmp;

r7_54_tmp <= r6[54];
r7[54] <= r7_54_tmp;

r7_55_tmp <= r6[55];
r7[55] <= r7_55_tmp;

r7_56_tmp <= r6[56];
r7[56] <= r7_56_tmp;

r7_57_tmp <= r6[57];
r7[57] <= r7_57_tmp;

r7_58_tmp <= r6[58];
r7[58] <= r7_58_tmp;

r7_59_tmp <= r6[59];
r7[59] <= r7_59_tmp;

r7_60_tmp <= r6[60];
r7[60] <= r7_60_tmp;

r7_61_tmp <= r6[61];
r7[61] <= r7_61_tmp;

r7_62_tmp <= r6[62];
r7[62] <= r7_62_tmp;

r7_63_tmp <= r6[63];
r7[63] <= r7_63_tmp;

r7_72_tmp <= r6[72];
r7[72] <= r7_72_tmp;

r7_73_tmp <= r6[73];
r7[73] <= r7_73_tmp;

r7_74_tmp <= r6[74];
r7[74] <= r7_74_tmp;

r7_75_tmp <= r6[75];
r7[75] <= r7_75_tmp;

r7_76_tmp <= r6[76];
r7[76] <= r7_76_tmp;

r7_77_tmp <= r6[77];
r7[77] <= r7_77_tmp;

r7_78_tmp <= r6[78];
r7[78] <= r7_78_tmp;

r7_79_tmp <= r6[79];
r7[79] <= r7_79_tmp;

//--------------------------
//---------layer : 8------------
cmp196_in0 <= r7[8];
cmp196_in1 <= r7[32];
r8[8] <= cmp196_out0;
r8[32] <= cmp196_out1;

cmp197_in0 <= r7[9];
cmp197_in1 <= r7[33];
r8[9] <= cmp197_out0;
r8[33] <= cmp197_out1;

cmp198_in0 <= r7[10];
cmp198_in1 <= r7[34];
r8[10] <= cmp198_out0;
r8[34] <= cmp198_out1;

cmp199_in0 <= r7[11];
cmp199_in1 <= r7[35];
r8[11] <= cmp199_out0;
r8[35] <= cmp199_out1;

cmp200_in0 <= r7[12];
cmp200_in1 <= r7[36];
r8[12] <= cmp200_out0;
r8[36] <= cmp200_out1;

cmp201_in0 <= r7[13];
cmp201_in1 <= r7[37];
r8[13] <= cmp201_out0;
r8[37] <= cmp201_out1;

cmp202_in0 <= r7[14];
cmp202_in1 <= r7[38];
r8[14] <= cmp202_out0;
r8[38] <= cmp202_out1;

cmp203_in0 <= r7[15];
cmp203_in1 <= r7[39];
r8[15] <= cmp203_out0;
r8[39] <= cmp203_out1;

cmp204_in0 <= r7[24];
cmp204_in1 <= r7[48];
r8[24] <= cmp204_out0;
r8[48] <= cmp204_out1;

cmp205_in0 <= r7[25];
cmp205_in1 <= r7[49];
r8[25] <= cmp205_out0;
r8[49] <= cmp205_out1;

cmp206_in0 <= r7[26];
cmp206_in1 <= r7[50];
r8[26] <= cmp206_out0;
r8[50] <= cmp206_out1;

cmp207_in0 <= r7[27];
cmp207_in1 <= r7[51];
r8[27] <= cmp207_out0;
r8[51] <= cmp207_out1;

cmp208_in0 <= r7[28];
cmp208_in1 <= r7[52];
r8[28] <= cmp208_out0;
r8[52] <= cmp208_out1;

cmp209_in0 <= r7[29];
cmp209_in1 <= r7[53];
r8[29] <= cmp209_out0;
r8[53] <= cmp209_out1;

cmp210_in0 <= r7[30];
cmp210_in1 <= r7[54];
r8[30] <= cmp210_out0;
r8[54] <= cmp210_out1;

cmp211_in0 <= r7[31];
cmp211_in1 <= r7[55];
r8[31] <= cmp211_out0;
r8[55] <= cmp211_out1;

cmp212_in0 <= r7[40];
cmp212_in1 <= r7[64];
r8[40] <= cmp212_out0;
r8[64] <= cmp212_out1;

cmp213_in0 <= r7[41];
cmp213_in1 <= r7[65];
r8[41] <= cmp213_out0;
r8[65] <= cmp213_out1;

cmp214_in0 <= r7[42];
cmp214_in1 <= r7[66];
r8[42] <= cmp214_out0;
r8[66] <= cmp214_out1;

cmp215_in0 <= r7[43];
cmp215_in1 <= r7[67];
r8[43] <= cmp215_out0;
r8[67] <= cmp215_out1;

cmp216_in0 <= r7[44];
cmp216_in1 <= r7[68];
r8[44] <= cmp216_out0;
r8[68] <= cmp216_out1;

cmp217_in0 <= r7[45];
cmp217_in1 <= r7[69];
r8[45] <= cmp217_out0;
r8[69] <= cmp217_out1;

cmp218_in0 <= r7[46];
cmp218_in1 <= r7[70];
r8[46] <= cmp218_out0;
r8[70] <= cmp218_out1;

cmp219_in0 <= r7[47];
cmp219_in1 <= r7[71];
r8[47] <= cmp219_out0;
r8[71] <= cmp219_out1;

cmp220_in0 <= r7[56];
cmp220_in1 <= r7[80];
r8[56] <= cmp220_out0;
r8[80] <= cmp220_out1;

r8_0_tmp <= r7[0];
r8[0] <= r8_0_tmp;

r8_1_tmp <= r7[1];
r8[1] <= r8_1_tmp;

r8_2_tmp <= r7[2];
r8[2] <= r8_2_tmp;

r8_3_tmp <= r7[3];
r8[3] <= r8_3_tmp;

r8_4_tmp <= r7[4];
r8[4] <= r8_4_tmp;

r8_5_tmp <= r7[5];
r8[5] <= r8_5_tmp;

r8_6_tmp <= r7[6];
r8[6] <= r8_6_tmp;

r8_7_tmp <= r7[7];
r8[7] <= r8_7_tmp;

r8_16_tmp <= r7[16];
r8[16] <= r8_16_tmp;

r8_17_tmp <= r7[17];
r8[17] <= r8_17_tmp;

r8_18_tmp <= r7[18];
r8[18] <= r8_18_tmp;

r8_19_tmp <= r7[19];
r8[19] <= r8_19_tmp;

r8_20_tmp <= r7[20];
r8[20] <= r8_20_tmp;

r8_21_tmp <= r7[21];
r8[21] <= r8_21_tmp;

r8_22_tmp <= r7[22];
r8[22] <= r8_22_tmp;

r8_23_tmp <= r7[23];
r8[23] <= r8_23_tmp;

r8_57_tmp <= r7[57];
r8[57] <= r8_57_tmp;

r8_58_tmp <= r7[58];
r8[58] <= r8_58_tmp;

r8_59_tmp <= r7[59];
r8[59] <= r8_59_tmp;

r8_60_tmp <= r7[60];
r8[60] <= r8_60_tmp;

r8_61_tmp <= r7[61];
r8[61] <= r8_61_tmp;

r8_62_tmp <= r7[62];
r8[62] <= r8_62_tmp;

r8_63_tmp <= r7[63];
r8[63] <= r8_63_tmp;

r8_72_tmp <= r7[72];
r8[72] <= r8_72_tmp;

r8_73_tmp <= r7[73];
r8[73] <= r8_73_tmp;

r8_74_tmp <= r7[74];
r8[74] <= r8_74_tmp;

r8_75_tmp <= r7[75];
r8[75] <= r8_75_tmp;

r8_76_tmp <= r7[76];
r8[76] <= r8_76_tmp;

r8_77_tmp <= r7[77];
r8[77] <= r8_77_tmp;

r8_78_tmp <= r7[78];
r8[78] <= r8_78_tmp;

r8_79_tmp <= r7[79];
r8[79] <= r8_79_tmp;

//--------------------------
//---------layer : 9------------
cmp221_in0 <= r8[8];
cmp221_in1 <= r8[16];
r9[8] <= cmp221_out0;
r9[16] <= cmp221_out1;

cmp222_in0 <= r8[9];
cmp222_in1 <= r8[17];
r9[9] <= cmp222_out0;
r9[17] <= cmp222_out1;

cmp223_in0 <= r8[10];
cmp223_in1 <= r8[18];
r9[10] <= cmp223_out0;
r9[18] <= cmp223_out1;

cmp224_in0 <= r8[11];
cmp224_in1 <= r8[19];
r9[11] <= cmp224_out0;
r9[19] <= cmp224_out1;

cmp225_in0 <= r8[12];
cmp225_in1 <= r8[20];
r9[12] <= cmp225_out0;
r9[20] <= cmp225_out1;

cmp226_in0 <= r8[13];
cmp226_in1 <= r8[21];
r9[13] <= cmp226_out0;
r9[21] <= cmp226_out1;

cmp227_in0 <= r8[14];
cmp227_in1 <= r8[22];
r9[14] <= cmp227_out0;
r9[22] <= cmp227_out1;

cmp228_in0 <= r8[15];
cmp228_in1 <= r8[23];
r9[15] <= cmp228_out0;
r9[23] <= cmp228_out1;

cmp229_in0 <= r8[24];
cmp229_in1 <= r8[32];
r9[24] <= cmp229_out0;
r9[32] <= cmp229_out1;

cmp230_in0 <= r8[25];
cmp230_in1 <= r8[33];
r9[25] <= cmp230_out0;
r9[33] <= cmp230_out1;

cmp231_in0 <= r8[26];
cmp231_in1 <= r8[34];
r9[26] <= cmp231_out0;
r9[34] <= cmp231_out1;

cmp232_in0 <= r8[27];
cmp232_in1 <= r8[35];
r9[27] <= cmp232_out0;
r9[35] <= cmp232_out1;

cmp233_in0 <= r8[28];
cmp233_in1 <= r8[36];
r9[28] <= cmp233_out0;
r9[36] <= cmp233_out1;

cmp234_in0 <= r8[29];
cmp234_in1 <= r8[37];
r9[29] <= cmp234_out0;
r9[37] <= cmp234_out1;

cmp235_in0 <= r8[30];
cmp235_in1 <= r8[38];
r9[30] <= cmp235_out0;
r9[38] <= cmp235_out1;

cmp236_in0 <= r8[31];
cmp236_in1 <= r8[39];
r9[31] <= cmp236_out0;
r9[39] <= cmp236_out1;

cmp237_in0 <= r8[40];
cmp237_in1 <= r8[48];
r9[40] <= cmp237_out0;
r9[48] <= cmp237_out1;

cmp238_in0 <= r8[41];
cmp238_in1 <= r8[49];
r9[41] <= cmp238_out0;
r9[49] <= cmp238_out1;

cmp239_in0 <= r8[42];
cmp239_in1 <= r8[50];
r9[42] <= cmp239_out0;
r9[50] <= cmp239_out1;

cmp240_in0 <= r8[43];
cmp240_in1 <= r8[51];
r9[43] <= cmp240_out0;
r9[51] <= cmp240_out1;

cmp241_in0 <= r8[44];
cmp241_in1 <= r8[52];
r9[44] <= cmp241_out0;
r9[52] <= cmp241_out1;

cmp242_in0 <= r8[45];
cmp242_in1 <= r8[53];
r9[45] <= cmp242_out0;
r9[53] <= cmp242_out1;

cmp243_in0 <= r8[46];
cmp243_in1 <= r8[54];
r9[46] <= cmp243_out0;
r9[54] <= cmp243_out1;

cmp244_in0 <= r8[47];
cmp244_in1 <= r8[55];
r9[47] <= cmp244_out0;
r9[55] <= cmp244_out1;

cmp245_in0 <= r8[56];
cmp245_in1 <= r8[64];
r9[56] <= cmp245_out0;
r9[64] <= cmp245_out1;

cmp246_in0 <= r8[57];
cmp246_in1 <= r8[65];
r9[57] <= cmp246_out0;
r9[65] <= cmp246_out1;

cmp247_in0 <= r8[58];
cmp247_in1 <= r8[66];
r9[58] <= cmp247_out0;
r9[66] <= cmp247_out1;

cmp248_in0 <= r8[59];
cmp248_in1 <= r8[67];
r9[59] <= cmp248_out0;
r9[67] <= cmp248_out1;

cmp249_in0 <= r8[60];
cmp249_in1 <= r8[68];
r9[60] <= cmp249_out0;
r9[68] <= cmp249_out1;

cmp250_in0 <= r8[61];
cmp250_in1 <= r8[69];
r9[61] <= cmp250_out0;
r9[69] <= cmp250_out1;

cmp251_in0 <= r8[62];
cmp251_in1 <= r8[70];
r9[62] <= cmp251_out0;
r9[70] <= cmp251_out1;

cmp252_in0 <= r8[63];
cmp252_in1 <= r8[71];
r9[63] <= cmp252_out0;
r9[71] <= cmp252_out1;

cmp253_in0 <= r8[72];
cmp253_in1 <= r8[80];
r9[72] <= cmp253_out0;
r9[80] <= cmp253_out1;

cmp254_in0 <= r8[0];
cmp254_in1 <= r8[4];
r9[0] <= cmp254_out0;
r9[4] <= cmp254_out1;

cmp255_in0 <= r8[1];
cmp255_in1 <= r8[5];
r9[1] <= cmp255_out0;
r9[5] <= cmp255_out1;

cmp256_in0 <= r8[2];
cmp256_in1 <= r8[6];
r9[2] <= cmp256_out0;
r9[6] <= cmp256_out1;

cmp257_in0 <= r8[3];
cmp257_in1 <= r8[7];
r9[3] <= cmp257_out0;
r9[7] <= cmp257_out1;

r9_73_tmp <= r8[73];
r9[73] <= r9_73_tmp;

r9_74_tmp <= r8[74];
r9[74] <= r9_74_tmp;

r9_75_tmp <= r8[75];
r9[75] <= r9_75_tmp;

r9_76_tmp <= r8[76];
r9[76] <= r9_76_tmp;

r9_77_tmp <= r8[77];
r9[77] <= r9_77_tmp;

r9_78_tmp <= r8[78];
r9[78] <= r9_78_tmp;

r9_79_tmp <= r8[79];
r9[79] <= r9_79_tmp;

//--------------------------
//---------layer : 10------------
cmp258_in0 <= r9[8];
cmp258_in1 <= r9[12];
r10[8] <= cmp258_out0;
r10[12] <= cmp258_out1;

cmp259_in0 <= r9[9];
cmp259_in1 <= r9[13];
r10[9] <= cmp259_out0;
r10[13] <= cmp259_out1;

cmp260_in0 <= r9[10];
cmp260_in1 <= r9[14];
r10[10] <= cmp260_out0;
r10[14] <= cmp260_out1;

cmp261_in0 <= r9[11];
cmp261_in1 <= r9[15];
r10[11] <= cmp261_out0;
r10[15] <= cmp261_out1;

cmp262_in0 <= r9[16];
cmp262_in1 <= r9[20];
r10[16] <= cmp262_out0;
r10[20] <= cmp262_out1;

cmp263_in0 <= r9[17];
cmp263_in1 <= r9[21];
r10[17] <= cmp263_out0;
r10[21] <= cmp263_out1;

cmp264_in0 <= r9[18];
cmp264_in1 <= r9[22];
r10[18] <= cmp264_out0;
r10[22] <= cmp264_out1;

cmp265_in0 <= r9[19];
cmp265_in1 <= r9[23];
r10[19] <= cmp265_out0;
r10[23] <= cmp265_out1;

cmp266_in0 <= r9[24];
cmp266_in1 <= r9[28];
r10[24] <= cmp266_out0;
r10[28] <= cmp266_out1;

cmp267_in0 <= r9[25];
cmp267_in1 <= r9[29];
r10[25] <= cmp267_out0;
r10[29] <= cmp267_out1;

cmp268_in0 <= r9[26];
cmp268_in1 <= r9[30];
r10[26] <= cmp268_out0;
r10[30] <= cmp268_out1;

cmp269_in0 <= r9[27];
cmp269_in1 <= r9[31];
r10[27] <= cmp269_out0;
r10[31] <= cmp269_out1;

cmp270_in0 <= r9[32];
cmp270_in1 <= r9[36];
r10[32] <= cmp270_out0;
r10[36] <= cmp270_out1;

cmp271_in0 <= r9[33];
cmp271_in1 <= r9[37];
r10[33] <= cmp271_out0;
r10[37] <= cmp271_out1;

cmp272_in0 <= r9[34];
cmp272_in1 <= r9[38];
r10[34] <= cmp272_out0;
r10[38] <= cmp272_out1;

cmp273_in0 <= r9[35];
cmp273_in1 <= r9[39];
r10[35] <= cmp273_out0;
r10[39] <= cmp273_out1;

cmp274_in0 <= r9[40];
cmp274_in1 <= r9[44];
r10[40] <= cmp274_out0;
r10[44] <= cmp274_out1;

cmp275_in0 <= r9[41];
cmp275_in1 <= r9[45];
r10[41] <= cmp275_out0;
r10[45] <= cmp275_out1;

cmp276_in0 <= r9[42];
cmp276_in1 <= r9[46];
r10[42] <= cmp276_out0;
r10[46] <= cmp276_out1;

cmp277_in0 <= r9[43];
cmp277_in1 <= r9[47];
r10[43] <= cmp277_out0;
r10[47] <= cmp277_out1;

cmp278_in0 <= r9[48];
cmp278_in1 <= r9[52];
r10[48] <= cmp278_out0;
r10[52] <= cmp278_out1;

cmp279_in0 <= r9[49];
cmp279_in1 <= r9[53];
r10[49] <= cmp279_out0;
r10[53] <= cmp279_out1;

cmp280_in0 <= r9[50];
cmp280_in1 <= r9[54];
r10[50] <= cmp280_out0;
r10[54] <= cmp280_out1;

cmp281_in0 <= r9[51];
cmp281_in1 <= r9[55];
r10[51] <= cmp281_out0;
r10[55] <= cmp281_out1;

cmp282_in0 <= r9[56];
cmp282_in1 <= r9[60];
r10[56] <= cmp282_out0;
r10[60] <= cmp282_out1;

cmp283_in0 <= r9[57];
cmp283_in1 <= r9[61];
r10[57] <= cmp283_out0;
r10[61] <= cmp283_out1;

cmp284_in0 <= r9[58];
cmp284_in1 <= r9[62];
r10[58] <= cmp284_out0;
r10[62] <= cmp284_out1;

cmp285_in0 <= r9[59];
cmp285_in1 <= r9[63];
r10[59] <= cmp285_out0;
r10[63] <= cmp285_out1;

cmp286_in0 <= r9[64];
cmp286_in1 <= r9[68];
r10[64] <= cmp286_out0;
r10[68] <= cmp286_out1;

cmp287_in0 <= r9[65];
cmp287_in1 <= r9[69];
r10[65] <= cmp287_out0;
r10[69] <= cmp287_out1;

cmp288_in0 <= r9[66];
cmp288_in1 <= r9[70];
r10[66] <= cmp288_out0;
r10[70] <= cmp288_out1;

cmp289_in0 <= r9[67];
cmp289_in1 <= r9[71];
r10[67] <= cmp289_out0;
r10[71] <= cmp289_out1;

cmp290_in0 <= r9[72];
cmp290_in1 <= r9[76];
r10[72] <= cmp290_out0;
r10[76] <= cmp290_out1;

cmp291_in0 <= r9[73];
cmp291_in1 <= r9[77];
r10[73] <= cmp291_out0;
r10[77] <= cmp291_out1;

cmp292_in0 <= r9[74];
cmp292_in1 <= r9[78];
r10[74] <= cmp292_out0;
r10[78] <= cmp292_out1;

cmp293_in0 <= r9[75];
cmp293_in1 <= r9[79];
r10[75] <= cmp293_out0;
r10[79] <= cmp293_out1;

r10_0_tmp <= r9[0];
r10[0] <= r10_0_tmp;

r10_1_tmp <= r9[1];
r10[1] <= r10_1_tmp;

r10_2_tmp <= r9[2];
r10[2] <= r10_2_tmp;

r10_3_tmp <= r9[3];
r10[3] <= r10_3_tmp;

r10_4_tmp <= r9[4];
r10[4] <= r10_4_tmp;

r10_5_tmp <= r9[5];
r10[5] <= r10_5_tmp;

r10_6_tmp <= r9[6];
r10[6] <= r10_6_tmp;

r10_7_tmp <= r9[7];
r10[7] <= r10_7_tmp;

r10_80_tmp <= r9[80];
r10[80] <= r10_80_tmp;

//--------------------------
//---------layer : 11------------
cmp294_in0 <= r10[4];
cmp294_in1 <= r10[64];
r11[4] <= cmp294_out0;
r11[64] <= cmp294_out1;

cmp295_in0 <= r10[5];
cmp295_in1 <= r10[65];
r11[5] <= cmp295_out0;
r11[65] <= cmp295_out1;

cmp296_in0 <= r10[6];
cmp296_in1 <= r10[66];
r11[6] <= cmp296_out0;
r11[66] <= cmp296_out1;

cmp297_in0 <= r10[7];
cmp297_in1 <= r10[67];
r11[7] <= cmp297_out0;
r11[67] <= cmp297_out1;

cmp298_in0 <= r10[12];
cmp298_in1 <= r10[72];
r11[12] <= cmp298_out0;
r11[72] <= cmp298_out1;

cmp299_in0 <= r10[13];
cmp299_in1 <= r10[73];
r11[13] <= cmp299_out0;
r11[73] <= cmp299_out1;

cmp300_in0 <= r10[14];
cmp300_in1 <= r10[74];
r11[14] <= cmp300_out0;
r11[74] <= cmp300_out1;

cmp301_in0 <= r10[15];
cmp301_in1 <= r10[75];
r11[15] <= cmp301_out0;
r11[75] <= cmp301_out1;

cmp302_in0 <= r10[20];
cmp302_in1 <= r10[80];
r11[20] <= cmp302_out0;
r11[80] <= cmp302_out1;

r11_0_tmp <= r10[0];
r11[0] <= r11_0_tmp;

r11_1_tmp <= r10[1];
r11[1] <= r11_1_tmp;

r11_2_tmp <= r10[2];
r11[2] <= r11_2_tmp;

r11_3_tmp <= r10[3];
r11[3] <= r11_3_tmp;

r11_8_tmp <= r10[8];
r11[8] <= r11_8_tmp;

r11_9_tmp <= r10[9];
r11[9] <= r11_9_tmp;

r11_10_tmp <= r10[10];
r11[10] <= r11_10_tmp;

r11_11_tmp <= r10[11];
r11[11] <= r11_11_tmp;

r11_16_tmp <= r10[16];
r11[16] <= r11_16_tmp;

r11_17_tmp <= r10[17];
r11[17] <= r11_17_tmp;

r11_18_tmp <= r10[18];
r11[18] <= r11_18_tmp;

r11_19_tmp <= r10[19];
r11[19] <= r11_19_tmp;

r11_21_tmp <= r10[21];
r11[21] <= r11_21_tmp;

r11_22_tmp <= r10[22];
r11[22] <= r11_22_tmp;

r11_23_tmp <= r10[23];
r11[23] <= r11_23_tmp;

r11_24_tmp <= r10[24];
r11[24] <= r11_24_tmp;

r11_25_tmp <= r10[25];
r11[25] <= r11_25_tmp;

r11_26_tmp <= r10[26];
r11[26] <= r11_26_tmp;

r11_27_tmp <= r10[27];
r11[27] <= r11_27_tmp;

r11_28_tmp <= r10[28];
r11[28] <= r11_28_tmp;

r11_29_tmp <= r10[29];
r11[29] <= r11_29_tmp;

r11_30_tmp <= r10[30];
r11[30] <= r11_30_tmp;

r11_31_tmp <= r10[31];
r11[31] <= r11_31_tmp;

r11_32_tmp <= r10[32];
r11[32] <= r11_32_tmp;

r11_33_tmp <= r10[33];
r11[33] <= r11_33_tmp;

r11_34_tmp <= r10[34];
r11[34] <= r11_34_tmp;

r11_35_tmp <= r10[35];
r11[35] <= r11_35_tmp;

r11_36_tmp <= r10[36];
r11[36] <= r11_36_tmp;

r11_37_tmp <= r10[37];
r11[37] <= r11_37_tmp;

r11_38_tmp <= r10[38];
r11[38] <= r11_38_tmp;

r11_39_tmp <= r10[39];
r11[39] <= r11_39_tmp;

r11_40_tmp <= r10[40];
r11[40] <= r11_40_tmp;

r11_41_tmp <= r10[41];
r11[41] <= r11_41_tmp;

r11_42_tmp <= r10[42];
r11[42] <= r11_42_tmp;

r11_43_tmp <= r10[43];
r11[43] <= r11_43_tmp;

r11_44_tmp <= r10[44];
r11[44] <= r11_44_tmp;

r11_45_tmp <= r10[45];
r11[45] <= r11_45_tmp;

r11_46_tmp <= r10[46];
r11[46] <= r11_46_tmp;

r11_47_tmp <= r10[47];
r11[47] <= r11_47_tmp;

r11_48_tmp <= r10[48];
r11[48] <= r11_48_tmp;

r11_49_tmp <= r10[49];
r11[49] <= r11_49_tmp;

r11_50_tmp <= r10[50];
r11[50] <= r11_50_tmp;

r11_51_tmp <= r10[51];
r11[51] <= r11_51_tmp;

r11_52_tmp <= r10[52];
r11[52] <= r11_52_tmp;

r11_53_tmp <= r10[53];
r11[53] <= r11_53_tmp;

r11_54_tmp <= r10[54];
r11[54] <= r11_54_tmp;

r11_55_tmp <= r10[55];
r11[55] <= r11_55_tmp;

r11_56_tmp <= r10[56];
r11[56] <= r11_56_tmp;

r11_57_tmp <= r10[57];
r11[57] <= r11_57_tmp;

r11_58_tmp <= r10[58];
r11[58] <= r11_58_tmp;

r11_59_tmp <= r10[59];
r11[59] <= r11_59_tmp;

r11_60_tmp <= r10[60];
r11[60] <= r11_60_tmp;

r11_61_tmp <= r10[61];
r11[61] <= r11_61_tmp;

r11_62_tmp <= r10[62];
r11[62] <= r11_62_tmp;

r11_63_tmp <= r10[63];
r11[63] <= r11_63_tmp;

r11_68_tmp <= r10[68];
r11[68] <= r11_68_tmp;

r11_69_tmp <= r10[69];
r11[69] <= r11_69_tmp;

r11_70_tmp <= r10[70];
r11[70] <= r11_70_tmp;

r11_71_tmp <= r10[71];
r11[71] <= r11_71_tmp;

r11_76_tmp <= r10[76];
r11[76] <= r11_76_tmp;

r11_77_tmp <= r10[77];
r11[77] <= r11_77_tmp;

r11_78_tmp <= r10[78];
r11[78] <= r11_78_tmp;

r11_79_tmp <= r10[79];
r11[79] <= r11_79_tmp;

//--------------------------
//---------layer : 12------------
cmp303_in0 <= r11[4];
cmp303_in1 <= r11[32];
r12[4] <= cmp303_out0;
r12[32] <= cmp303_out1;

cmp304_in0 <= r11[5];
cmp304_in1 <= r11[33];
r12[5] <= cmp304_out0;
r12[33] <= cmp304_out1;

cmp305_in0 <= r11[6];
cmp305_in1 <= r11[34];
r12[6] <= cmp305_out0;
r12[34] <= cmp305_out1;

cmp306_in0 <= r11[7];
cmp306_in1 <= r11[35];
r12[7] <= cmp306_out0;
r12[35] <= cmp306_out1;

cmp307_in0 <= r11[12];
cmp307_in1 <= r11[40];
r12[12] <= cmp307_out0;
r12[40] <= cmp307_out1;

cmp308_in0 <= r11[13];
cmp308_in1 <= r11[41];
r12[13] <= cmp308_out0;
r12[41] <= cmp308_out1;

cmp309_in0 <= r11[14];
cmp309_in1 <= r11[42];
r12[14] <= cmp309_out0;
r12[42] <= cmp309_out1;

cmp310_in0 <= r11[15];
cmp310_in1 <= r11[43];
r12[15] <= cmp310_out0;
r12[43] <= cmp310_out1;

cmp311_in0 <= r11[20];
cmp311_in1 <= r11[48];
r12[20] <= cmp311_out0;
r12[48] <= cmp311_out1;

cmp312_in0 <= r11[21];
cmp312_in1 <= r11[49];
r12[21] <= cmp312_out0;
r12[49] <= cmp312_out1;

cmp313_in0 <= r11[22];
cmp313_in1 <= r11[50];
r12[22] <= cmp313_out0;
r12[50] <= cmp313_out1;

cmp314_in0 <= r11[23];
cmp314_in1 <= r11[51];
r12[23] <= cmp314_out0;
r12[51] <= cmp314_out1;

cmp315_in0 <= r11[28];
cmp315_in1 <= r11[56];
r12[28] <= cmp315_out0;
r12[56] <= cmp315_out1;

cmp316_in0 <= r11[29];
cmp316_in1 <= r11[57];
r12[29] <= cmp316_out0;
r12[57] <= cmp316_out1;

cmp317_in0 <= r11[30];
cmp317_in1 <= r11[58];
r12[30] <= cmp317_out0;
r12[58] <= cmp317_out1;

cmp318_in0 <= r11[31];
cmp318_in1 <= r11[59];
r12[31] <= cmp318_out0;
r12[59] <= cmp318_out1;

cmp319_in0 <= r11[36];
cmp319_in1 <= r11[64];
r12[36] <= cmp319_out0;
r12[64] <= cmp319_out1;

cmp320_in0 <= r11[37];
cmp320_in1 <= r11[65];
r12[37] <= cmp320_out0;
r12[65] <= cmp320_out1;

cmp321_in0 <= r11[38];
cmp321_in1 <= r11[66];
r12[38] <= cmp321_out0;
r12[66] <= cmp321_out1;

cmp322_in0 <= r11[39];
cmp322_in1 <= r11[67];
r12[39] <= cmp322_out0;
r12[67] <= cmp322_out1;

cmp323_in0 <= r11[44];
cmp323_in1 <= r11[72];
r12[44] <= cmp323_out0;
r12[72] <= cmp323_out1;

cmp324_in0 <= r11[45];
cmp324_in1 <= r11[73];
r12[45] <= cmp324_out0;
r12[73] <= cmp324_out1;

cmp325_in0 <= r11[46];
cmp325_in1 <= r11[74];
r12[46] <= cmp325_out0;
r12[74] <= cmp325_out1;

cmp326_in0 <= r11[47];
cmp326_in1 <= r11[75];
r12[47] <= cmp326_out0;
r12[75] <= cmp326_out1;

cmp327_in0 <= r11[52];
cmp327_in1 <= r11[80];
r12[52] <= cmp327_out0;
r12[80] <= cmp327_out1;

r12_0_tmp <= r11[0];
r12[0] <= r12_0_tmp;

r12_1_tmp <= r11[1];
r12[1] <= r12_1_tmp;

r12_2_tmp <= r11[2];
r12[2] <= r12_2_tmp;

r12_3_tmp <= r11[3];
r12[3] <= r12_3_tmp;

r12_8_tmp <= r11[8];
r12[8] <= r12_8_tmp;

r12_9_tmp <= r11[9];
r12[9] <= r12_9_tmp;

r12_10_tmp <= r11[10];
r12[10] <= r12_10_tmp;

r12_11_tmp <= r11[11];
r12[11] <= r12_11_tmp;

r12_16_tmp <= r11[16];
r12[16] <= r12_16_tmp;

r12_17_tmp <= r11[17];
r12[17] <= r12_17_tmp;

r12_18_tmp <= r11[18];
r12[18] <= r12_18_tmp;

r12_19_tmp <= r11[19];
r12[19] <= r12_19_tmp;

r12_24_tmp <= r11[24];
r12[24] <= r12_24_tmp;

r12_25_tmp <= r11[25];
r12[25] <= r12_25_tmp;

r12_26_tmp <= r11[26];
r12[26] <= r12_26_tmp;

r12_27_tmp <= r11[27];
r12[27] <= r12_27_tmp;

r12_53_tmp <= r11[53];
r12[53] <= r12_53_tmp;

r12_54_tmp <= r11[54];
r12[54] <= r12_54_tmp;

r12_55_tmp <= r11[55];
r12[55] <= r12_55_tmp;

r12_60_tmp <= r11[60];
r12[60] <= r12_60_tmp;

r12_61_tmp <= r11[61];
r12[61] <= r12_61_tmp;

r12_62_tmp <= r11[62];
r12[62] <= r12_62_tmp;

r12_63_tmp <= r11[63];
r12[63] <= r12_63_tmp;

r12_68_tmp <= r11[68];
r12[68] <= r12_68_tmp;

r12_69_tmp <= r11[69];
r12[69] <= r12_69_tmp;

r12_70_tmp <= r11[70];
r12[70] <= r12_70_tmp;

r12_71_tmp <= r11[71];
r12[71] <= r12_71_tmp;

r12_76_tmp <= r11[76];
r12[76] <= r12_76_tmp;

r12_77_tmp <= r11[77];
r12[77] <= r12_77_tmp;

r12_78_tmp <= r11[78];
r12[78] <= r12_78_tmp;

r12_79_tmp <= r11[79];
r12[79] <= r12_79_tmp;

//--------------------------
//---------layer : 13------------
cmp328_in0 <= r12[4];
cmp328_in1 <= r12[16];
r13[4] <= cmp328_out0;
r13[16] <= cmp328_out1;

cmp329_in0 <= r12[5];
cmp329_in1 <= r12[17];
r13[5] <= cmp329_out0;
r13[17] <= cmp329_out1;

cmp330_in0 <= r12[6];
cmp330_in1 <= r12[18];
r13[6] <= cmp330_out0;
r13[18] <= cmp330_out1;

cmp331_in0 <= r12[7];
cmp331_in1 <= r12[19];
r13[7] <= cmp331_out0;
r13[19] <= cmp331_out1;

cmp332_in0 <= r12[12];
cmp332_in1 <= r12[24];
r13[12] <= cmp332_out0;
r13[24] <= cmp332_out1;

cmp333_in0 <= r12[13];
cmp333_in1 <= r12[25];
r13[13] <= cmp333_out0;
r13[25] <= cmp333_out1;

cmp334_in0 <= r12[14];
cmp334_in1 <= r12[26];
r13[14] <= cmp334_out0;
r13[26] <= cmp334_out1;

cmp335_in0 <= r12[15];
cmp335_in1 <= r12[27];
r13[15] <= cmp335_out0;
r13[27] <= cmp335_out1;

cmp336_in0 <= r12[20];
cmp336_in1 <= r12[32];
r13[20] <= cmp336_out0;
r13[32] <= cmp336_out1;

cmp337_in0 <= r12[21];
cmp337_in1 <= r12[33];
r13[21] <= cmp337_out0;
r13[33] <= cmp337_out1;

cmp338_in0 <= r12[22];
cmp338_in1 <= r12[34];
r13[22] <= cmp338_out0;
r13[34] <= cmp338_out1;

cmp339_in0 <= r12[23];
cmp339_in1 <= r12[35];
r13[23] <= cmp339_out0;
r13[35] <= cmp339_out1;

cmp340_in0 <= r12[28];
cmp340_in1 <= r12[40];
r13[28] <= cmp340_out0;
r13[40] <= cmp340_out1;

cmp341_in0 <= r12[29];
cmp341_in1 <= r12[41];
r13[29] <= cmp341_out0;
r13[41] <= cmp341_out1;

cmp342_in0 <= r12[30];
cmp342_in1 <= r12[42];
r13[30] <= cmp342_out0;
r13[42] <= cmp342_out1;

cmp343_in0 <= r12[31];
cmp343_in1 <= r12[43];
r13[31] <= cmp343_out0;
r13[43] <= cmp343_out1;

cmp344_in0 <= r12[36];
cmp344_in1 <= r12[48];
r13[36] <= cmp344_out0;
r13[48] <= cmp344_out1;

cmp345_in0 <= r12[37];
cmp345_in1 <= r12[49];
r13[37] <= cmp345_out0;
r13[49] <= cmp345_out1;

cmp346_in0 <= r12[38];
cmp346_in1 <= r12[50];
r13[38] <= cmp346_out0;
r13[50] <= cmp346_out1;

cmp347_in0 <= r12[39];
cmp347_in1 <= r12[51];
r13[39] <= cmp347_out0;
r13[51] <= cmp347_out1;

cmp348_in0 <= r12[44];
cmp348_in1 <= r12[56];
r13[44] <= cmp348_out0;
r13[56] <= cmp348_out1;

cmp349_in0 <= r12[45];
cmp349_in1 <= r12[57];
r13[45] <= cmp349_out0;
r13[57] <= cmp349_out1;

cmp350_in0 <= r12[46];
cmp350_in1 <= r12[58];
r13[46] <= cmp350_out0;
r13[58] <= cmp350_out1;

cmp351_in0 <= r12[47];
cmp351_in1 <= r12[59];
r13[47] <= cmp351_out0;
r13[59] <= cmp351_out1;

cmp352_in0 <= r12[52];
cmp352_in1 <= r12[64];
r13[52] <= cmp352_out0;
r13[64] <= cmp352_out1;

cmp353_in0 <= r12[53];
cmp353_in1 <= r12[65];
r13[53] <= cmp353_out0;
r13[65] <= cmp353_out1;

cmp354_in0 <= r12[54];
cmp354_in1 <= r12[66];
r13[54] <= cmp354_out0;
r13[66] <= cmp354_out1;

cmp355_in0 <= r12[55];
cmp355_in1 <= r12[67];
r13[55] <= cmp355_out0;
r13[67] <= cmp355_out1;

cmp356_in0 <= r12[60];
cmp356_in1 <= r12[72];
r13[60] <= cmp356_out0;
r13[72] <= cmp356_out1;

cmp357_in0 <= r12[61];
cmp357_in1 <= r12[73];
r13[61] <= cmp357_out0;
r13[73] <= cmp357_out1;

cmp358_in0 <= r12[62];
cmp358_in1 <= r12[74];
r13[62] <= cmp358_out0;
r13[74] <= cmp358_out1;

cmp359_in0 <= r12[63];
cmp359_in1 <= r12[75];
r13[63] <= cmp359_out0;
r13[75] <= cmp359_out1;

cmp360_in0 <= r12[68];
cmp360_in1 <= r12[80];
r13[68] <= cmp360_out0;
r13[80] <= cmp360_out1;

r13_0_tmp <= r12[0];
r13[0] <= r13_0_tmp;

r13_1_tmp <= r12[1];
r13[1] <= r13_1_tmp;

r13_2_tmp <= r12[2];
r13[2] <= r13_2_tmp;

r13_3_tmp <= r12[3];
r13[3] <= r13_3_tmp;

r13_8_tmp <= r12[8];
r13[8] <= r13_8_tmp;

r13_9_tmp <= r12[9];
r13[9] <= r13_9_tmp;

r13_10_tmp <= r12[10];
r13[10] <= r13_10_tmp;

r13_11_tmp <= r12[11];
r13[11] <= r13_11_tmp;

r13_69_tmp <= r12[69];
r13[69] <= r13_69_tmp;

r13_70_tmp <= r12[70];
r13[70] <= r13_70_tmp;

r13_71_tmp <= r12[71];
r13[71] <= r13_71_tmp;

r13_76_tmp <= r12[76];
r13[76] <= r13_76_tmp;

r13_77_tmp <= r12[77];
r13[77] <= r13_77_tmp;

r13_78_tmp <= r12[78];
r13[78] <= r13_78_tmp;

r13_79_tmp <= r12[79];
r13[79] <= r13_79_tmp;

//--------------------------
//---------layer : 14------------
cmp361_in0 <= r13[4];
cmp361_in1 <= r13[8];
r14[4] <= cmp361_out0;
r14[8] <= cmp361_out1;

cmp362_in0 <= r13[5];
cmp362_in1 <= r13[9];
r14[5] <= cmp362_out0;
r14[9] <= cmp362_out1;

cmp363_in0 <= r13[6];
cmp363_in1 <= r13[10];
r14[6] <= cmp363_out0;
r14[10] <= cmp363_out1;

cmp364_in0 <= r13[7];
cmp364_in1 <= r13[11];
r14[7] <= cmp364_out0;
r14[11] <= cmp364_out1;

cmp365_in0 <= r13[12];
cmp365_in1 <= r13[16];
r14[12] <= cmp365_out0;
r14[16] <= cmp365_out1;

cmp366_in0 <= r13[13];
cmp366_in1 <= r13[17];
r14[13] <= cmp366_out0;
r14[17] <= cmp366_out1;

cmp367_in0 <= r13[14];
cmp367_in1 <= r13[18];
r14[14] <= cmp367_out0;
r14[18] <= cmp367_out1;

cmp368_in0 <= r13[15];
cmp368_in1 <= r13[19];
r14[15] <= cmp368_out0;
r14[19] <= cmp368_out1;

cmp369_in0 <= r13[20];
cmp369_in1 <= r13[24];
r14[20] <= cmp369_out0;
r14[24] <= cmp369_out1;

cmp370_in0 <= r13[21];
cmp370_in1 <= r13[25];
r14[21] <= cmp370_out0;
r14[25] <= cmp370_out1;

cmp371_in0 <= r13[22];
cmp371_in1 <= r13[26];
r14[22] <= cmp371_out0;
r14[26] <= cmp371_out1;

cmp372_in0 <= r13[23];
cmp372_in1 <= r13[27];
r14[23] <= cmp372_out0;
r14[27] <= cmp372_out1;

cmp373_in0 <= r13[28];
cmp373_in1 <= r13[32];
r14[28] <= cmp373_out0;
r14[32] <= cmp373_out1;

cmp374_in0 <= r13[29];
cmp374_in1 <= r13[33];
r14[29] <= cmp374_out0;
r14[33] <= cmp374_out1;

cmp375_in0 <= r13[30];
cmp375_in1 <= r13[34];
r14[30] <= cmp375_out0;
r14[34] <= cmp375_out1;

cmp376_in0 <= r13[31];
cmp376_in1 <= r13[35];
r14[31] <= cmp376_out0;
r14[35] <= cmp376_out1;

cmp377_in0 <= r13[36];
cmp377_in1 <= r13[40];
r14[36] <= cmp377_out0;
r14[40] <= cmp377_out1;

cmp378_in0 <= r13[37];
cmp378_in1 <= r13[41];
r14[37] <= cmp378_out0;
r14[41] <= cmp378_out1;

cmp379_in0 <= r13[38];
cmp379_in1 <= r13[42];
r14[38] <= cmp379_out0;
r14[42] <= cmp379_out1;

cmp380_in0 <= r13[39];
cmp380_in1 <= r13[43];
r14[39] <= cmp380_out0;
r14[43] <= cmp380_out1;

cmp381_in0 <= r13[44];
cmp381_in1 <= r13[48];
r14[44] <= cmp381_out0;
r14[48] <= cmp381_out1;

cmp382_in0 <= r13[45];
cmp382_in1 <= r13[49];
r14[45] <= cmp382_out0;
r14[49] <= cmp382_out1;

cmp383_in0 <= r13[46];
cmp383_in1 <= r13[50];
r14[46] <= cmp383_out0;
r14[50] <= cmp383_out1;

cmp384_in0 <= r13[47];
cmp384_in1 <= r13[51];
r14[47] <= cmp384_out0;
r14[51] <= cmp384_out1;

cmp385_in0 <= r13[52];
cmp385_in1 <= r13[56];
r14[52] <= cmp385_out0;
r14[56] <= cmp385_out1;

cmp386_in0 <= r13[53];
cmp386_in1 <= r13[57];
r14[53] <= cmp386_out0;
r14[57] <= cmp386_out1;

cmp387_in0 <= r13[54];
cmp387_in1 <= r13[58];
r14[54] <= cmp387_out0;
r14[58] <= cmp387_out1;

cmp388_in0 <= r13[55];
cmp388_in1 <= r13[59];
r14[55] <= cmp388_out0;
r14[59] <= cmp388_out1;

cmp389_in0 <= r13[60];
cmp389_in1 <= r13[64];
r14[60] <= cmp389_out0;
r14[64] <= cmp389_out1;

cmp390_in0 <= r13[61];
cmp390_in1 <= r13[65];
r14[61] <= cmp390_out0;
r14[65] <= cmp390_out1;

cmp391_in0 <= r13[62];
cmp391_in1 <= r13[66];
r14[62] <= cmp391_out0;
r14[66] <= cmp391_out1;

cmp392_in0 <= r13[63];
cmp392_in1 <= r13[67];
r14[63] <= cmp392_out0;
r14[67] <= cmp392_out1;

cmp393_in0 <= r13[68];
cmp393_in1 <= r13[72];
r14[68] <= cmp393_out0;
r14[72] <= cmp393_out1;

cmp394_in0 <= r13[69];
cmp394_in1 <= r13[73];
r14[69] <= cmp394_out0;
r14[73] <= cmp394_out1;

cmp395_in0 <= r13[70];
cmp395_in1 <= r13[74];
r14[70] <= cmp395_out0;
r14[74] <= cmp395_out1;

cmp396_in0 <= r13[71];
cmp396_in1 <= r13[75];
r14[71] <= cmp396_out0;
r14[75] <= cmp396_out1;

cmp397_in0 <= r13[76];
cmp397_in1 <= r13[80];
r14[76] <= cmp397_out0;
r14[80] <= cmp397_out1;

cmp398_in0 <= r13[0];
cmp398_in1 <= r13[2];
r14[0] <= cmp398_out0;
r14[2] <= cmp398_out1;

cmp399_in0 <= r13[1];
cmp399_in1 <= r13[3];
r14[1] <= cmp399_out0;
r14[3] <= cmp399_out1;

r14_77_tmp <= r13[77];
r14[77] <= r14_77_tmp;

r14_78_tmp <= r13[78];
r14[78] <= r14_78_tmp;

r14_79_tmp <= r13[79];
r14[79] <= r14_79_tmp;

//--------------------------
//---------layer : 15------------
cmp400_in0 <= r14[4];
cmp400_in1 <= r14[6];
r15[4] <= cmp400_out0;
r15[6] <= cmp400_out1;

cmp401_in0 <= r14[5];
cmp401_in1 <= r14[7];
r15[5] <= cmp401_out0;
r15[7] <= cmp401_out1;

cmp402_in0 <= r14[8];
cmp402_in1 <= r14[10];
r15[8] <= cmp402_out0;
r15[10] <= cmp402_out1;

cmp403_in0 <= r14[9];
cmp403_in1 <= r14[11];
r15[9] <= cmp403_out0;
r15[11] <= cmp403_out1;

cmp404_in0 <= r14[12];
cmp404_in1 <= r14[14];
r15[12] <= cmp404_out0;
r15[14] <= cmp404_out1;

cmp405_in0 <= r14[13];
cmp405_in1 <= r14[15];
r15[13] <= cmp405_out0;
r15[15] <= cmp405_out1;

cmp406_in0 <= r14[16];
cmp406_in1 <= r14[18];
r15[16] <= cmp406_out0;
r15[18] <= cmp406_out1;

cmp407_in0 <= r14[17];
cmp407_in1 <= r14[19];
r15[17] <= cmp407_out0;
r15[19] <= cmp407_out1;

cmp408_in0 <= r14[20];
cmp408_in1 <= r14[22];
r15[20] <= cmp408_out0;
r15[22] <= cmp408_out1;

cmp409_in0 <= r14[21];
cmp409_in1 <= r14[23];
r15[21] <= cmp409_out0;
r15[23] <= cmp409_out1;

cmp410_in0 <= r14[24];
cmp410_in1 <= r14[26];
r15[24] <= cmp410_out0;
r15[26] <= cmp410_out1;

cmp411_in0 <= r14[25];
cmp411_in1 <= r14[27];
r15[25] <= cmp411_out0;
r15[27] <= cmp411_out1;

cmp412_in0 <= r14[28];
cmp412_in1 <= r14[30];
r15[28] <= cmp412_out0;
r15[30] <= cmp412_out1;

cmp413_in0 <= r14[29];
cmp413_in1 <= r14[31];
r15[29] <= cmp413_out0;
r15[31] <= cmp413_out1;

cmp414_in0 <= r14[32];
cmp414_in1 <= r14[34];
r15[32] <= cmp414_out0;
r15[34] <= cmp414_out1;

cmp415_in0 <= r14[33];
cmp415_in1 <= r14[35];
r15[33] <= cmp415_out0;
r15[35] <= cmp415_out1;

cmp416_in0 <= r14[36];
cmp416_in1 <= r14[38];
r15[36] <= cmp416_out0;
r15[38] <= cmp416_out1;

cmp417_in0 <= r14[37];
cmp417_in1 <= r14[39];
r15[37] <= cmp417_out0;
r15[39] <= cmp417_out1;

cmp418_in0 <= r14[40];
cmp418_in1 <= r14[42];
r15[40] <= cmp418_out0;
r15[42] <= cmp418_out1;

cmp419_in0 <= r14[41];
cmp419_in1 <= r14[43];
r15[41] <= cmp419_out0;
r15[43] <= cmp419_out1;

cmp420_in0 <= r14[44];
cmp420_in1 <= r14[46];
r15[44] <= cmp420_out0;
r15[46] <= cmp420_out1;

cmp421_in0 <= r14[45];
cmp421_in1 <= r14[47];
r15[45] <= cmp421_out0;
r15[47] <= cmp421_out1;

cmp422_in0 <= r14[48];
cmp422_in1 <= r14[50];
r15[48] <= cmp422_out0;
r15[50] <= cmp422_out1;

cmp423_in0 <= r14[49];
cmp423_in1 <= r14[51];
r15[49] <= cmp423_out0;
r15[51] <= cmp423_out1;

cmp424_in0 <= r14[52];
cmp424_in1 <= r14[54];
r15[52] <= cmp424_out0;
r15[54] <= cmp424_out1;

cmp425_in0 <= r14[53];
cmp425_in1 <= r14[55];
r15[53] <= cmp425_out0;
r15[55] <= cmp425_out1;

cmp426_in0 <= r14[56];
cmp426_in1 <= r14[58];
r15[56] <= cmp426_out0;
r15[58] <= cmp426_out1;

cmp427_in0 <= r14[57];
cmp427_in1 <= r14[59];
r15[57] <= cmp427_out0;
r15[59] <= cmp427_out1;

cmp428_in0 <= r14[60];
cmp428_in1 <= r14[62];
r15[60] <= cmp428_out0;
r15[62] <= cmp428_out1;

cmp429_in0 <= r14[61];
cmp429_in1 <= r14[63];
r15[61] <= cmp429_out0;
r15[63] <= cmp429_out1;

cmp430_in0 <= r14[64];
cmp430_in1 <= r14[66];
r15[64] <= cmp430_out0;
r15[66] <= cmp430_out1;

cmp431_in0 <= r14[65];
cmp431_in1 <= r14[67];
r15[65] <= cmp431_out0;
r15[67] <= cmp431_out1;

cmp432_in0 <= r14[68];
cmp432_in1 <= r14[70];
r15[68] <= cmp432_out0;
r15[70] <= cmp432_out1;

cmp433_in0 <= r14[69];
cmp433_in1 <= r14[71];
r15[69] <= cmp433_out0;
r15[71] <= cmp433_out1;

cmp434_in0 <= r14[72];
cmp434_in1 <= r14[74];
r15[72] <= cmp434_out0;
r15[74] <= cmp434_out1;

cmp435_in0 <= r14[73];
cmp435_in1 <= r14[75];
r15[73] <= cmp435_out0;
r15[75] <= cmp435_out1;

cmp436_in0 <= r14[76];
cmp436_in1 <= r14[78];
r15[76] <= cmp436_out0;
r15[78] <= cmp436_out1;

cmp437_in0 <= r14[77];
cmp437_in1 <= r14[79];
r15[77] <= cmp437_out0;
r15[79] <= cmp437_out1;

r15_0_tmp <= r14[0];
r15[0] <= r15_0_tmp;

r15_1_tmp <= r14[1];
r15[1] <= r15_1_tmp;

r15_2_tmp <= r14[2];
r15[2] <= r15_2_tmp;

r15_3_tmp <= r14[3];
r15[3] <= r15_3_tmp;

r15_80_tmp <= r14[80];
r15[80] <= r15_80_tmp;

//--------------------------
//---------layer : 16------------
cmp438_in0 <= r15[2];
cmp438_in1 <= r15[64];
r16[2] <= cmp438_out0;
r16[64] <= cmp438_out1;

cmp439_in0 <= r15[3];
cmp439_in1 <= r15[65];
r16[3] <= cmp439_out0;
r16[65] <= cmp439_out1;

cmp440_in0 <= r15[6];
cmp440_in1 <= r15[68];
r16[6] <= cmp440_out0;
r16[68] <= cmp440_out1;

cmp441_in0 <= r15[7];
cmp441_in1 <= r15[69];
r16[7] <= cmp441_out0;
r16[69] <= cmp441_out1;

cmp442_in0 <= r15[10];
cmp442_in1 <= r15[72];
r16[10] <= cmp442_out0;
r16[72] <= cmp442_out1;

cmp443_in0 <= r15[11];
cmp443_in1 <= r15[73];
r16[11] <= cmp443_out0;
r16[73] <= cmp443_out1;

cmp444_in0 <= r15[14];
cmp444_in1 <= r15[76];
r16[14] <= cmp444_out0;
r16[76] <= cmp444_out1;

cmp445_in0 <= r15[15];
cmp445_in1 <= r15[77];
r16[15] <= cmp445_out0;
r16[77] <= cmp445_out1;

cmp446_in0 <= r15[18];
cmp446_in1 <= r15[80];
r16[18] <= cmp446_out0;
r16[80] <= cmp446_out1;

r16_0_tmp <= r15[0];
r16[0] <= r16_0_tmp;

r16_1_tmp <= r15[1];
r16[1] <= r16_1_tmp;

r16_4_tmp <= r15[4];
r16[4] <= r16_4_tmp;

r16_5_tmp <= r15[5];
r16[5] <= r16_5_tmp;

r16_8_tmp <= r15[8];
r16[8] <= r16_8_tmp;

r16_9_tmp <= r15[9];
r16[9] <= r16_9_tmp;

r16_12_tmp <= r15[12];
r16[12] <= r16_12_tmp;

r16_13_tmp <= r15[13];
r16[13] <= r16_13_tmp;

r16_16_tmp <= r15[16];
r16[16] <= r16_16_tmp;

r16_17_tmp <= r15[17];
r16[17] <= r16_17_tmp;

r16_19_tmp <= r15[19];
r16[19] <= r16_19_tmp;

r16_20_tmp <= r15[20];
r16[20] <= r16_20_tmp;

r16_21_tmp <= r15[21];
r16[21] <= r16_21_tmp;

r16_22_tmp <= r15[22];
r16[22] <= r16_22_tmp;

r16_23_tmp <= r15[23];
r16[23] <= r16_23_tmp;

r16_24_tmp <= r15[24];
r16[24] <= r16_24_tmp;

r16_25_tmp <= r15[25];
r16[25] <= r16_25_tmp;

r16_26_tmp <= r15[26];
r16[26] <= r16_26_tmp;

r16_27_tmp <= r15[27];
r16[27] <= r16_27_tmp;

r16_28_tmp <= r15[28];
r16[28] <= r16_28_tmp;

r16_29_tmp <= r15[29];
r16[29] <= r16_29_tmp;

r16_30_tmp <= r15[30];
r16[30] <= r16_30_tmp;

r16_31_tmp <= r15[31];
r16[31] <= r16_31_tmp;

r16_32_tmp <= r15[32];
r16[32] <= r16_32_tmp;

r16_33_tmp <= r15[33];
r16[33] <= r16_33_tmp;

r16_34_tmp <= r15[34];
r16[34] <= r16_34_tmp;

r16_35_tmp <= r15[35];
r16[35] <= r16_35_tmp;

r16_36_tmp <= r15[36];
r16[36] <= r16_36_tmp;

r16_37_tmp <= r15[37];
r16[37] <= r16_37_tmp;

r16_38_tmp <= r15[38];
r16[38] <= r16_38_tmp;

r16_39_tmp <= r15[39];
r16[39] <= r16_39_tmp;

r16_40_tmp <= r15[40];
r16[40] <= r16_40_tmp;

r16_41_tmp <= r15[41];
r16[41] <= r16_41_tmp;

r16_42_tmp <= r15[42];
r16[42] <= r16_42_tmp;

r16_43_tmp <= r15[43];
r16[43] <= r16_43_tmp;

r16_44_tmp <= r15[44];
r16[44] <= r16_44_tmp;

r16_45_tmp <= r15[45];
r16[45] <= r16_45_tmp;

r16_46_tmp <= r15[46];
r16[46] <= r16_46_tmp;

r16_47_tmp <= r15[47];
r16[47] <= r16_47_tmp;

r16_48_tmp <= r15[48];
r16[48] <= r16_48_tmp;

r16_49_tmp <= r15[49];
r16[49] <= r16_49_tmp;

r16_50_tmp <= r15[50];
r16[50] <= r16_50_tmp;

r16_51_tmp <= r15[51];
r16[51] <= r16_51_tmp;

r16_52_tmp <= r15[52];
r16[52] <= r16_52_tmp;

r16_53_tmp <= r15[53];
r16[53] <= r16_53_tmp;

r16_54_tmp <= r15[54];
r16[54] <= r16_54_tmp;

r16_55_tmp <= r15[55];
r16[55] <= r16_55_tmp;

r16_56_tmp <= r15[56];
r16[56] <= r16_56_tmp;

r16_57_tmp <= r15[57];
r16[57] <= r16_57_tmp;

r16_58_tmp <= r15[58];
r16[58] <= r16_58_tmp;

r16_59_tmp <= r15[59];
r16[59] <= r16_59_tmp;

r16_60_tmp <= r15[60];
r16[60] <= r16_60_tmp;

r16_61_tmp <= r15[61];
r16[61] <= r16_61_tmp;

r16_62_tmp <= r15[62];
r16[62] <= r16_62_tmp;

r16_63_tmp <= r15[63];
r16[63] <= r16_63_tmp;

r16_66_tmp <= r15[66];
r16[66] <= r16_66_tmp;

r16_67_tmp <= r15[67];
r16[67] <= r16_67_tmp;

r16_70_tmp <= r15[70];
r16[70] <= r16_70_tmp;

r16_71_tmp <= r15[71];
r16[71] <= r16_71_tmp;

r16_74_tmp <= r15[74];
r16[74] <= r16_74_tmp;

r16_75_tmp <= r15[75];
r16[75] <= r16_75_tmp;

r16_78_tmp <= r15[78];
r16[78] <= r16_78_tmp;

r16_79_tmp <= r15[79];
r16[79] <= r16_79_tmp;

//--------------------------
//---------layer : 17------------
cmp447_in0 <= r16[2];
cmp447_in1 <= r16[32];
r17[2] <= cmp447_out0;
r17[32] <= cmp447_out1;

cmp448_in0 <= r16[3];
cmp448_in1 <= r16[33];
r17[3] <= cmp448_out0;
r17[33] <= cmp448_out1;

cmp449_in0 <= r16[6];
cmp449_in1 <= r16[36];
r17[6] <= cmp449_out0;
r17[36] <= cmp449_out1;

cmp450_in0 <= r16[7];
cmp450_in1 <= r16[37];
r17[7] <= cmp450_out0;
r17[37] <= cmp450_out1;

cmp451_in0 <= r16[10];
cmp451_in1 <= r16[40];
r17[10] <= cmp451_out0;
r17[40] <= cmp451_out1;

cmp452_in0 <= r16[11];
cmp452_in1 <= r16[41];
r17[11] <= cmp452_out0;
r17[41] <= cmp452_out1;

cmp453_in0 <= r16[14];
cmp453_in1 <= r16[44];
r17[14] <= cmp453_out0;
r17[44] <= cmp453_out1;

cmp454_in0 <= r16[15];
cmp454_in1 <= r16[45];
r17[15] <= cmp454_out0;
r17[45] <= cmp454_out1;

cmp455_in0 <= r16[18];
cmp455_in1 <= r16[48];
r17[18] <= cmp455_out0;
r17[48] <= cmp455_out1;

cmp456_in0 <= r16[19];
cmp456_in1 <= r16[49];
r17[19] <= cmp456_out0;
r17[49] <= cmp456_out1;

cmp457_in0 <= r16[22];
cmp457_in1 <= r16[52];
r17[22] <= cmp457_out0;
r17[52] <= cmp457_out1;

cmp458_in0 <= r16[23];
cmp458_in1 <= r16[53];
r17[23] <= cmp458_out0;
r17[53] <= cmp458_out1;

cmp459_in0 <= r16[26];
cmp459_in1 <= r16[56];
r17[26] <= cmp459_out0;
r17[56] <= cmp459_out1;

cmp460_in0 <= r16[27];
cmp460_in1 <= r16[57];
r17[27] <= cmp460_out0;
r17[57] <= cmp460_out1;

cmp461_in0 <= r16[30];
cmp461_in1 <= r16[60];
r17[30] <= cmp461_out0;
r17[60] <= cmp461_out1;

cmp462_in0 <= r16[31];
cmp462_in1 <= r16[61];
r17[31] <= cmp462_out0;
r17[61] <= cmp462_out1;

cmp463_in0 <= r16[34];
cmp463_in1 <= r16[64];
r17[34] <= cmp463_out0;
r17[64] <= cmp463_out1;

cmp464_in0 <= r16[35];
cmp464_in1 <= r16[65];
r17[35] <= cmp464_out0;
r17[65] <= cmp464_out1;

cmp465_in0 <= r16[38];
cmp465_in1 <= r16[68];
r17[38] <= cmp465_out0;
r17[68] <= cmp465_out1;

cmp466_in0 <= r16[39];
cmp466_in1 <= r16[69];
r17[39] <= cmp466_out0;
r17[69] <= cmp466_out1;

cmp467_in0 <= r16[42];
cmp467_in1 <= r16[72];
r17[42] <= cmp467_out0;
r17[72] <= cmp467_out1;

cmp468_in0 <= r16[43];
cmp468_in1 <= r16[73];
r17[43] <= cmp468_out0;
r17[73] <= cmp468_out1;

cmp469_in0 <= r16[46];
cmp469_in1 <= r16[76];
r17[46] <= cmp469_out0;
r17[76] <= cmp469_out1;

cmp470_in0 <= r16[47];
cmp470_in1 <= r16[77];
r17[47] <= cmp470_out0;
r17[77] <= cmp470_out1;

cmp471_in0 <= r16[50];
cmp471_in1 <= r16[80];
r17[50] <= cmp471_out0;
r17[80] <= cmp471_out1;

r17_0_tmp <= r16[0];
r17[0] <= r17_0_tmp;

r17_1_tmp <= r16[1];
r17[1] <= r17_1_tmp;

r17_4_tmp <= r16[4];
r17[4] <= r17_4_tmp;

r17_5_tmp <= r16[5];
r17[5] <= r17_5_tmp;

r17_8_tmp <= r16[8];
r17[8] <= r17_8_tmp;

r17_9_tmp <= r16[9];
r17[9] <= r17_9_tmp;

r17_12_tmp <= r16[12];
r17[12] <= r17_12_tmp;

r17_13_tmp <= r16[13];
r17[13] <= r17_13_tmp;

r17_16_tmp <= r16[16];
r17[16] <= r17_16_tmp;

r17_17_tmp <= r16[17];
r17[17] <= r17_17_tmp;

r17_20_tmp <= r16[20];
r17[20] <= r17_20_tmp;

r17_21_tmp <= r16[21];
r17[21] <= r17_21_tmp;

r17_24_tmp <= r16[24];
r17[24] <= r17_24_tmp;

r17_25_tmp <= r16[25];
r17[25] <= r17_25_tmp;

r17_28_tmp <= r16[28];
r17[28] <= r17_28_tmp;

r17_29_tmp <= r16[29];
r17[29] <= r17_29_tmp;

r17_51_tmp <= r16[51];
r17[51] <= r17_51_tmp;

r17_54_tmp <= r16[54];
r17[54] <= r17_54_tmp;

r17_55_tmp <= r16[55];
r17[55] <= r17_55_tmp;

r17_58_tmp <= r16[58];
r17[58] <= r17_58_tmp;

r17_59_tmp <= r16[59];
r17[59] <= r17_59_tmp;

r17_62_tmp <= r16[62];
r17[62] <= r17_62_tmp;

r17_63_tmp <= r16[63];
r17[63] <= r17_63_tmp;

r17_66_tmp <= r16[66];
r17[66] <= r17_66_tmp;

r17_67_tmp <= r16[67];
r17[67] <= r17_67_tmp;

r17_70_tmp <= r16[70];
r17[70] <= r17_70_tmp;

r17_71_tmp <= r16[71];
r17[71] <= r17_71_tmp;

r17_74_tmp <= r16[74];
r17[74] <= r17_74_tmp;

r17_75_tmp <= r16[75];
r17[75] <= r17_75_tmp;

r17_78_tmp <= r16[78];
r17[78] <= r17_78_tmp;

r17_79_tmp <= r16[79];
r17[79] <= r17_79_tmp;

//--------------------------
//---------layer : 18------------
cmp472_in0 <= r17[2];
cmp472_in1 <= r17[16];
r18[2] <= cmp472_out0;
r18[16] <= cmp472_out1;

cmp473_in0 <= r17[3];
cmp473_in1 <= r17[17];
r18[3] <= cmp473_out0;
r18[17] <= cmp473_out1;

cmp474_in0 <= r17[6];
cmp474_in1 <= r17[20];
r18[6] <= cmp474_out0;
r18[20] <= cmp474_out1;

cmp475_in0 <= r17[7];
cmp475_in1 <= r17[21];
r18[7] <= cmp475_out0;
r18[21] <= cmp475_out1;

cmp476_in0 <= r17[10];
cmp476_in1 <= r17[24];
r18[10] <= cmp476_out0;
r18[24] <= cmp476_out1;

cmp477_in0 <= r17[11];
cmp477_in1 <= r17[25];
r18[11] <= cmp477_out0;
r18[25] <= cmp477_out1;

cmp478_in0 <= r17[14];
cmp478_in1 <= r17[28];
r18[14] <= cmp478_out0;
r18[28] <= cmp478_out1;

cmp479_in0 <= r17[15];
cmp479_in1 <= r17[29];
r18[15] <= cmp479_out0;
r18[29] <= cmp479_out1;

cmp480_in0 <= r17[18];
cmp480_in1 <= r17[32];
r18[18] <= cmp480_out0;
r18[32] <= cmp480_out1;

cmp481_in0 <= r17[19];
cmp481_in1 <= r17[33];
r18[19] <= cmp481_out0;
r18[33] <= cmp481_out1;

cmp482_in0 <= r17[22];
cmp482_in1 <= r17[36];
r18[22] <= cmp482_out0;
r18[36] <= cmp482_out1;

cmp483_in0 <= r17[23];
cmp483_in1 <= r17[37];
r18[23] <= cmp483_out0;
r18[37] <= cmp483_out1;

cmp484_in0 <= r17[26];
cmp484_in1 <= r17[40];
r18[26] <= cmp484_out0;
r18[40] <= cmp484_out1;

cmp485_in0 <= r17[27];
cmp485_in1 <= r17[41];
r18[27] <= cmp485_out0;
r18[41] <= cmp485_out1;

cmp486_in0 <= r17[30];
cmp486_in1 <= r17[44];
r18[30] <= cmp486_out0;
r18[44] <= cmp486_out1;

cmp487_in0 <= r17[31];
cmp487_in1 <= r17[45];
r18[31] <= cmp487_out0;
r18[45] <= cmp487_out1;

cmp488_in0 <= r17[34];
cmp488_in1 <= r17[48];
r18[34] <= cmp488_out0;
r18[48] <= cmp488_out1;

cmp489_in0 <= r17[35];
cmp489_in1 <= r17[49];
r18[35] <= cmp489_out0;
r18[49] <= cmp489_out1;

cmp490_in0 <= r17[38];
cmp490_in1 <= r17[52];
r18[38] <= cmp490_out0;
r18[52] <= cmp490_out1;

cmp491_in0 <= r17[39];
cmp491_in1 <= r17[53];
r18[39] <= cmp491_out0;
r18[53] <= cmp491_out1;

cmp492_in0 <= r17[42];
cmp492_in1 <= r17[56];
r18[42] <= cmp492_out0;
r18[56] <= cmp492_out1;

cmp493_in0 <= r17[43];
cmp493_in1 <= r17[57];
r18[43] <= cmp493_out0;
r18[57] <= cmp493_out1;

cmp494_in0 <= r17[46];
cmp494_in1 <= r17[60];
r18[46] <= cmp494_out0;
r18[60] <= cmp494_out1;

cmp495_in0 <= r17[47];
cmp495_in1 <= r17[61];
r18[47] <= cmp495_out0;
r18[61] <= cmp495_out1;

cmp496_in0 <= r17[50];
cmp496_in1 <= r17[64];
r18[50] <= cmp496_out0;
r18[64] <= cmp496_out1;

cmp497_in0 <= r17[51];
cmp497_in1 <= r17[65];
r18[51] <= cmp497_out0;
r18[65] <= cmp497_out1;

cmp498_in0 <= r17[54];
cmp498_in1 <= r17[68];
r18[54] <= cmp498_out0;
r18[68] <= cmp498_out1;

cmp499_in0 <= r17[55];
cmp499_in1 <= r17[69];
r18[55] <= cmp499_out0;
r18[69] <= cmp499_out1;

cmp500_in0 <= r17[58];
cmp500_in1 <= r17[72];
r18[58] <= cmp500_out0;
r18[72] <= cmp500_out1;

cmp501_in0 <= r17[59];
cmp501_in1 <= r17[73];
r18[59] <= cmp501_out0;
r18[73] <= cmp501_out1;

cmp502_in0 <= r17[62];
cmp502_in1 <= r17[76];
r18[62] <= cmp502_out0;
r18[76] <= cmp502_out1;

cmp503_in0 <= r17[63];
cmp503_in1 <= r17[77];
r18[63] <= cmp503_out0;
r18[77] <= cmp503_out1;

cmp504_in0 <= r17[66];
cmp504_in1 <= r17[80];
r18[66] <= cmp504_out0;
r18[80] <= cmp504_out1;

r18_0_tmp <= r17[0];
r18[0] <= r18_0_tmp;

r18_1_tmp <= r17[1];
r18[1] <= r18_1_tmp;

r18_4_tmp <= r17[4];
r18[4] <= r18_4_tmp;

r18_5_tmp <= r17[5];
r18[5] <= r18_5_tmp;

r18_8_tmp <= r17[8];
r18[8] <= r18_8_tmp;

r18_9_tmp <= r17[9];
r18[9] <= r18_9_tmp;

r18_12_tmp <= r17[12];
r18[12] <= r18_12_tmp;

r18_13_tmp <= r17[13];
r18[13] <= r18_13_tmp;

r18_67_tmp <= r17[67];
r18[67] <= r18_67_tmp;

r18_70_tmp <= r17[70];
r18[70] <= r18_70_tmp;

r18_71_tmp <= r17[71];
r18[71] <= r18_71_tmp;

r18_74_tmp <= r17[74];
r18[74] <= r18_74_tmp;

r18_75_tmp <= r17[75];
r18[75] <= r18_75_tmp;

r18_78_tmp <= r17[78];
r18[78] <= r18_78_tmp;

r18_79_tmp <= r17[79];
r18[79] <= r18_79_tmp;

//--------------------------
//---------layer : 19------------
cmp505_in0 <= r18[2];
cmp505_in1 <= r18[8];
r19[2] <= cmp505_out0;
r19[8] <= cmp505_out1;

cmp506_in0 <= r18[3];
cmp506_in1 <= r18[9];
r19[3] <= cmp506_out0;
r19[9] <= cmp506_out1;

cmp507_in0 <= r18[6];
cmp507_in1 <= r18[12];
r19[6] <= cmp507_out0;
r19[12] <= cmp507_out1;

cmp508_in0 <= r18[7];
cmp508_in1 <= r18[13];
r19[7] <= cmp508_out0;
r19[13] <= cmp508_out1;

cmp509_in0 <= r18[10];
cmp509_in1 <= r18[16];
r19[10] <= cmp509_out0;
r19[16] <= cmp509_out1;

cmp510_in0 <= r18[11];
cmp510_in1 <= r18[17];
r19[11] <= cmp510_out0;
r19[17] <= cmp510_out1;

cmp511_in0 <= r18[14];
cmp511_in1 <= r18[20];
r19[14] <= cmp511_out0;
r19[20] <= cmp511_out1;

cmp512_in0 <= r18[15];
cmp512_in1 <= r18[21];
r19[15] <= cmp512_out0;
r19[21] <= cmp512_out1;

cmp513_in0 <= r18[18];
cmp513_in1 <= r18[24];
r19[18] <= cmp513_out0;
r19[24] <= cmp513_out1;

cmp514_in0 <= r18[19];
cmp514_in1 <= r18[25];
r19[19] <= cmp514_out0;
r19[25] <= cmp514_out1;

cmp515_in0 <= r18[22];
cmp515_in1 <= r18[28];
r19[22] <= cmp515_out0;
r19[28] <= cmp515_out1;

cmp516_in0 <= r18[23];
cmp516_in1 <= r18[29];
r19[23] <= cmp516_out0;
r19[29] <= cmp516_out1;

cmp517_in0 <= r18[26];
cmp517_in1 <= r18[32];
r19[26] <= cmp517_out0;
r19[32] <= cmp517_out1;

cmp518_in0 <= r18[27];
cmp518_in1 <= r18[33];
r19[27] <= cmp518_out0;
r19[33] <= cmp518_out1;

cmp519_in0 <= r18[30];
cmp519_in1 <= r18[36];
r19[30] <= cmp519_out0;
r19[36] <= cmp519_out1;

cmp520_in0 <= r18[31];
cmp520_in1 <= r18[37];
r19[31] <= cmp520_out0;
r19[37] <= cmp520_out1;

cmp521_in0 <= r18[34];
cmp521_in1 <= r18[40];
r19[34] <= cmp521_out0;
r19[40] <= cmp521_out1;

cmp522_in0 <= r18[35];
cmp522_in1 <= r18[41];
r19[35] <= cmp522_out0;
r19[41] <= cmp522_out1;

cmp523_in0 <= r18[38];
cmp523_in1 <= r18[44];
r19[38] <= cmp523_out0;
r19[44] <= cmp523_out1;

cmp524_in0 <= r18[39];
cmp524_in1 <= r18[45];
r19[39] <= cmp524_out0;
r19[45] <= cmp524_out1;

cmp525_in0 <= r18[42];
cmp525_in1 <= r18[48];
r19[42] <= cmp525_out0;
r19[48] <= cmp525_out1;

cmp526_in0 <= r18[43];
cmp526_in1 <= r18[49];
r19[43] <= cmp526_out0;
r19[49] <= cmp526_out1;

cmp527_in0 <= r18[46];
cmp527_in1 <= r18[52];
r19[46] <= cmp527_out0;
r19[52] <= cmp527_out1;

cmp528_in0 <= r18[47];
cmp528_in1 <= r18[53];
r19[47] <= cmp528_out0;
r19[53] <= cmp528_out1;

cmp529_in0 <= r18[50];
cmp529_in1 <= r18[56];
r19[50] <= cmp529_out0;
r19[56] <= cmp529_out1;

cmp530_in0 <= r18[51];
cmp530_in1 <= r18[57];
r19[51] <= cmp530_out0;
r19[57] <= cmp530_out1;

cmp531_in0 <= r18[54];
cmp531_in1 <= r18[60];
r19[54] <= cmp531_out0;
r19[60] <= cmp531_out1;

cmp532_in0 <= r18[55];
cmp532_in1 <= r18[61];
r19[55] <= cmp532_out0;
r19[61] <= cmp532_out1;

cmp533_in0 <= r18[58];
cmp533_in1 <= r18[64];
r19[58] <= cmp533_out0;
r19[64] <= cmp533_out1;

cmp534_in0 <= r18[59];
cmp534_in1 <= r18[65];
r19[59] <= cmp534_out0;
r19[65] <= cmp534_out1;

cmp535_in0 <= r18[62];
cmp535_in1 <= r18[68];
r19[62] <= cmp535_out0;
r19[68] <= cmp535_out1;

cmp536_in0 <= r18[63];
cmp536_in1 <= r18[69];
r19[63] <= cmp536_out0;
r19[69] <= cmp536_out1;

cmp537_in0 <= r18[66];
cmp537_in1 <= r18[72];
r19[66] <= cmp537_out0;
r19[72] <= cmp537_out1;

cmp538_in0 <= r18[67];
cmp538_in1 <= r18[73];
r19[67] <= cmp538_out0;
r19[73] <= cmp538_out1;

cmp539_in0 <= r18[70];
cmp539_in1 <= r18[76];
r19[70] <= cmp539_out0;
r19[76] <= cmp539_out1;

cmp540_in0 <= r18[71];
cmp540_in1 <= r18[77];
r19[71] <= cmp540_out0;
r19[77] <= cmp540_out1;

cmp541_in0 <= r18[74];
cmp541_in1 <= r18[80];
r19[74] <= cmp541_out0;
r19[80] <= cmp541_out1;

r19_0_tmp <= r18[0];
r19[0] <= r19_0_tmp;

r19_1_tmp <= r18[1];
r19[1] <= r19_1_tmp;

r19_4_tmp <= r18[4];
r19[4] <= r19_4_tmp;

r19_5_tmp <= r18[5];
r19[5] <= r19_5_tmp;

r19_75_tmp <= r18[75];
r19[75] <= r19_75_tmp;

r19_78_tmp <= r18[78];
r19[78] <= r19_78_tmp;

r19_79_tmp <= r18[79];
r19[79] <= r19_79_tmp;

//--------------------------
//---------layer : 20------------
cmp542_in0 <= r19[2];
cmp542_in1 <= r19[4];
r20[2] <= cmp542_out0;
r20[4] <= cmp542_out1;

cmp543_in0 <= r19[3];
cmp543_in1 <= r19[5];
r20[3] <= cmp543_out0;
r20[5] <= cmp543_out1;

cmp544_in0 <= r19[6];
cmp544_in1 <= r19[8];
r20[6] <= cmp544_out0;
r20[8] <= cmp544_out1;

cmp545_in0 <= r19[7];
cmp545_in1 <= r19[9];
r20[7] <= cmp545_out0;
r20[9] <= cmp545_out1;

cmp546_in0 <= r19[10];
cmp546_in1 <= r19[12];
r20[10] <= cmp546_out0;
r20[12] <= cmp546_out1;

cmp547_in0 <= r19[11];
cmp547_in1 <= r19[13];
r20[11] <= cmp547_out0;
r20[13] <= cmp547_out1;

cmp548_in0 <= r19[14];
cmp548_in1 <= r19[16];
r20[14] <= cmp548_out0;
r20[16] <= cmp548_out1;

cmp549_in0 <= r19[15];
cmp549_in1 <= r19[17];
r20[15] <= cmp549_out0;
r20[17] <= cmp549_out1;

cmp550_in0 <= r19[18];
cmp550_in1 <= r19[20];
r20[18] <= cmp550_out0;
r20[20] <= cmp550_out1;

cmp551_in0 <= r19[19];
cmp551_in1 <= r19[21];
r20[19] <= cmp551_out0;
r20[21] <= cmp551_out1;

cmp552_in0 <= r19[22];
cmp552_in1 <= r19[24];
r20[22] <= cmp552_out0;
r20[24] <= cmp552_out1;

cmp553_in0 <= r19[23];
cmp553_in1 <= r19[25];
r20[23] <= cmp553_out0;
r20[25] <= cmp553_out1;

cmp554_in0 <= r19[26];
cmp554_in1 <= r19[28];
r20[26] <= cmp554_out0;
r20[28] <= cmp554_out1;

cmp555_in0 <= r19[27];
cmp555_in1 <= r19[29];
r20[27] <= cmp555_out0;
r20[29] <= cmp555_out1;

cmp556_in0 <= r19[30];
cmp556_in1 <= r19[32];
r20[30] <= cmp556_out0;
r20[32] <= cmp556_out1;

cmp557_in0 <= r19[31];
cmp557_in1 <= r19[33];
r20[31] <= cmp557_out0;
r20[33] <= cmp557_out1;

cmp558_in0 <= r19[34];
cmp558_in1 <= r19[36];
r20[34] <= cmp558_out0;
r20[36] <= cmp558_out1;

cmp559_in0 <= r19[35];
cmp559_in1 <= r19[37];
r20[35] <= cmp559_out0;
r20[37] <= cmp559_out1;

cmp560_in0 <= r19[38];
cmp560_in1 <= r19[40];
r20[38] <= cmp560_out0;
r20[40] <= cmp560_out1;

cmp561_in0 <= r19[39];
cmp561_in1 <= r19[41];
r20[39] <= cmp561_out0;
r20[41] <= cmp561_out1;

cmp562_in0 <= r19[42];
cmp562_in1 <= r19[44];
r20[42] <= cmp562_out0;
r20[44] <= cmp562_out1;

cmp563_in0 <= r19[43];
cmp563_in1 <= r19[45];
r20[43] <= cmp563_out0;
r20[45] <= cmp563_out1;

cmp564_in0 <= r19[46];
cmp564_in1 <= r19[48];
r20[46] <= cmp564_out0;
r20[48] <= cmp564_out1;

cmp565_in0 <= r19[47];
cmp565_in1 <= r19[49];
r20[47] <= cmp565_out0;
r20[49] <= cmp565_out1;

cmp566_in0 <= r19[50];
cmp566_in1 <= r19[52];
r20[50] <= cmp566_out0;
r20[52] <= cmp566_out1;

cmp567_in0 <= r19[51];
cmp567_in1 <= r19[53];
r20[51] <= cmp567_out0;
r20[53] <= cmp567_out1;

cmp568_in0 <= r19[54];
cmp568_in1 <= r19[56];
r20[54] <= cmp568_out0;
r20[56] <= cmp568_out1;

cmp569_in0 <= r19[55];
cmp569_in1 <= r19[57];
r20[55] <= cmp569_out0;
r20[57] <= cmp569_out1;

cmp570_in0 <= r19[58];
cmp570_in1 <= r19[60];
r20[58] <= cmp570_out0;
r20[60] <= cmp570_out1;

cmp571_in0 <= r19[59];
cmp571_in1 <= r19[61];
r20[59] <= cmp571_out0;
r20[61] <= cmp571_out1;

cmp572_in0 <= r19[62];
cmp572_in1 <= r19[64];
r20[62] <= cmp572_out0;
r20[64] <= cmp572_out1;

cmp573_in0 <= r19[63];
cmp573_in1 <= r19[65];
r20[63] <= cmp573_out0;
r20[65] <= cmp573_out1;

cmp574_in0 <= r19[66];
cmp574_in1 <= r19[68];
r20[66] <= cmp574_out0;
r20[68] <= cmp574_out1;

cmp575_in0 <= r19[67];
cmp575_in1 <= r19[69];
r20[67] <= cmp575_out0;
r20[69] <= cmp575_out1;

cmp576_in0 <= r19[70];
cmp576_in1 <= r19[72];
r20[70] <= cmp576_out0;
r20[72] <= cmp576_out1;

cmp577_in0 <= r19[71];
cmp577_in1 <= r19[73];
r20[71] <= cmp577_out0;
r20[73] <= cmp577_out1;

cmp578_in0 <= r19[74];
cmp578_in1 <= r19[76];
r20[74] <= cmp578_out0;
r20[76] <= cmp578_out1;

cmp579_in0 <= r19[75];
cmp579_in1 <= r19[77];
r20[75] <= cmp579_out0;
r20[77] <= cmp579_out1;

cmp580_in0 <= r19[78];
cmp580_in1 <= r19[80];
r20[78] <= cmp580_out0;
r20[80] <= cmp580_out1;

cmp581_in0 <= r19[0];
cmp581_in1 <= r19[1];
r20[0] <= cmp581_out0;
r20[1] <= cmp581_out1;

r20_79_tmp <= r19[79];
r20[79] <= r20_79_tmp;

//--------------------------
//---------layer : 21------------
cmp582_in0 <= r20[2];
cmp582_in1 <= r20[3];
r21[2] <= cmp582_out0;
r21[3] <= cmp582_out1;

cmp583_in0 <= r20[4];
cmp583_in1 <= r20[5];
r21[4] <= cmp583_out0;
r21[5] <= cmp583_out1;

cmp584_in0 <= r20[6];
cmp584_in1 <= r20[7];
r21[6] <= cmp584_out0;
r21[7] <= cmp584_out1;

cmp585_in0 <= r20[8];
cmp585_in1 <= r20[9];
r21[8] <= cmp585_out0;
r21[9] <= cmp585_out1;

cmp586_in0 <= r20[10];
cmp586_in1 <= r20[11];
r21[10] <= cmp586_out0;
r21[11] <= cmp586_out1;

cmp587_in0 <= r20[12];
cmp587_in1 <= r20[13];
r21[12] <= cmp587_out0;
r21[13] <= cmp587_out1;

cmp588_in0 <= r20[14];
cmp588_in1 <= r20[15];
r21[14] <= cmp588_out0;
r21[15] <= cmp588_out1;

cmp589_in0 <= r20[16];
cmp589_in1 <= r20[17];
r21[16] <= cmp589_out0;
r21[17] <= cmp589_out1;

cmp590_in0 <= r20[18];
cmp590_in1 <= r20[19];
r21[18] <= cmp590_out0;
r21[19] <= cmp590_out1;

cmp591_in0 <= r20[20];
cmp591_in1 <= r20[21];
r21[20] <= cmp591_out0;
r21[21] <= cmp591_out1;

cmp592_in0 <= r20[22];
cmp592_in1 <= r20[23];
r21[22] <= cmp592_out0;
r21[23] <= cmp592_out1;

cmp593_in0 <= r20[24];
cmp593_in1 <= r20[25];
r21[24] <= cmp593_out0;
r21[25] <= cmp593_out1;

cmp594_in0 <= r20[26];
cmp594_in1 <= r20[27];
r21[26] <= cmp594_out0;
r21[27] <= cmp594_out1;

cmp595_in0 <= r20[28];
cmp595_in1 <= r20[29];
r21[28] <= cmp595_out0;
r21[29] <= cmp595_out1;

cmp596_in0 <= r20[30];
cmp596_in1 <= r20[31];
r21[30] <= cmp596_out0;
r21[31] <= cmp596_out1;

cmp597_in0 <= r20[32];
cmp597_in1 <= r20[33];
r21[32] <= cmp597_out0;
r21[33] <= cmp597_out1;

cmp598_in0 <= r20[34];
cmp598_in1 <= r20[35];
r21[34] <= cmp598_out0;
r21[35] <= cmp598_out1;

cmp599_in0 <= r20[36];
cmp599_in1 <= r20[37];
r21[36] <= cmp599_out0;
r21[37] <= cmp599_out1;

cmp600_in0 <= r20[38];
cmp600_in1 <= r20[39];
r21[38] <= cmp600_out0;
r21[39] <= cmp600_out1;

cmp601_in0 <= r20[40];
cmp601_in1 <= r20[41];
r21[40] <= cmp601_out0;
r21[41] <= cmp601_out1;

cmp602_in0 <= r20[42];
cmp602_in1 <= r20[43];
r21[42] <= cmp602_out0;
r21[43] <= cmp602_out1;

cmp603_in0 <= r20[44];
cmp603_in1 <= r20[45];
r21[44] <= cmp603_out0;
r21[45] <= cmp603_out1;

cmp604_in0 <= r20[46];
cmp604_in1 <= r20[47];
r21[46] <= cmp604_out0;
r21[47] <= cmp604_out1;

cmp605_in0 <= r20[48];
cmp605_in1 <= r20[49];
r21[48] <= cmp605_out0;
r21[49] <= cmp605_out1;

cmp606_in0 <= r20[50];
cmp606_in1 <= r20[51];
r21[50] <= cmp606_out0;
r21[51] <= cmp606_out1;

cmp607_in0 <= r20[52];
cmp607_in1 <= r20[53];
r21[52] <= cmp607_out0;
r21[53] <= cmp607_out1;

cmp608_in0 <= r20[54];
cmp608_in1 <= r20[55];
r21[54] <= cmp608_out0;
r21[55] <= cmp608_out1;

cmp609_in0 <= r20[56];
cmp609_in1 <= r20[57];
r21[56] <= cmp609_out0;
r21[57] <= cmp609_out1;

cmp610_in0 <= r20[58];
cmp610_in1 <= r20[59];
r21[58] <= cmp610_out0;
r21[59] <= cmp610_out1;

cmp611_in0 <= r20[60];
cmp611_in1 <= r20[61];
r21[60] <= cmp611_out0;
r21[61] <= cmp611_out1;

cmp612_in0 <= r20[62];
cmp612_in1 <= r20[63];
r21[62] <= cmp612_out0;
r21[63] <= cmp612_out1;

cmp613_in0 <= r20[64];
cmp613_in1 <= r20[65];
r21[64] <= cmp613_out0;
r21[65] <= cmp613_out1;

cmp614_in0 <= r20[66];
cmp614_in1 <= r20[67];
r21[66] <= cmp614_out0;
r21[67] <= cmp614_out1;

cmp615_in0 <= r20[68];
cmp615_in1 <= r20[69];
r21[68] <= cmp615_out0;
r21[69] <= cmp615_out1;

cmp616_in0 <= r20[70];
cmp616_in1 <= r20[71];
r21[70] <= cmp616_out0;
r21[71] <= cmp616_out1;

cmp617_in0 <= r20[72];
cmp617_in1 <= r20[73];
r21[72] <= cmp617_out0;
r21[73] <= cmp617_out1;

cmp618_in0 <= r20[74];
cmp618_in1 <= r20[75];
r21[74] <= cmp618_out0;
r21[75] <= cmp618_out1;

cmp619_in0 <= r20[76];
cmp619_in1 <= r20[77];
r21[76] <= cmp619_out0;
r21[77] <= cmp619_out1;

cmp620_in0 <= r20[78];
cmp620_in1 <= r20[79];
r21[78] <= cmp620_out0;
r21[79] <= cmp620_out1;

r21_0_tmp <= r20[0];
r21[0] <= r21_0_tmp;

r21_1_tmp <= r20[1];
r21[1] <= r21_1_tmp;

r21_80_tmp <= r20[80];
r21[80] <= r21_80_tmp;

//--------------------------
//---------layer : 22------------
cmp621_in0 <= r21[1];
cmp621_in1 <= r21[64];
r22[1] <= cmp621_out0;
r22[64] <= cmp621_out1;

cmp622_in0 <= r21[3];
cmp622_in1 <= r21[66];
r22[3] <= cmp622_out0;
r22[66] <= cmp622_out1;

cmp623_in0 <= r21[5];
cmp623_in1 <= r21[68];
r22[5] <= cmp623_out0;
r22[68] <= cmp623_out1;

cmp624_in0 <= r21[7];
cmp624_in1 <= r21[70];
r22[7] <= cmp624_out0;
r22[70] <= cmp624_out1;

cmp625_in0 <= r21[9];
cmp625_in1 <= r21[72];
r22[9] <= cmp625_out0;
r22[72] <= cmp625_out1;

cmp626_in0 <= r21[11];
cmp626_in1 <= r21[74];
r22[11] <= cmp626_out0;
r22[74] <= cmp626_out1;

cmp627_in0 <= r21[13];
cmp627_in1 <= r21[76];
r22[13] <= cmp627_out0;
r22[76] <= cmp627_out1;

cmp628_in0 <= r21[15];
cmp628_in1 <= r21[78];
r22[15] <= cmp628_out0;
r22[78] <= cmp628_out1;

cmp629_in0 <= r21[17];
cmp629_in1 <= r21[80];
r22[17] <= cmp629_out0;
r22[80] <= cmp629_out1;

r22_0_tmp <= r21[0];
r22[0] <= r22_0_tmp;

r22_2_tmp <= r21[2];
r22[2] <= r22_2_tmp;

r22_4_tmp <= r21[4];
r22[4] <= r22_4_tmp;

r22_6_tmp <= r21[6];
r22[6] <= r22_6_tmp;

r22_8_tmp <= r21[8];
r22[8] <= r22_8_tmp;

r22_10_tmp <= r21[10];
r22[10] <= r22_10_tmp;

r22_12_tmp <= r21[12];
r22[12] <= r22_12_tmp;

r22_14_tmp <= r21[14];
r22[14] <= r22_14_tmp;

r22_16_tmp <= r21[16];
r22[16] <= r22_16_tmp;

r22_18_tmp <= r21[18];
r22[18] <= r22_18_tmp;

r22_19_tmp <= r21[19];
r22[19] <= r22_19_tmp;

r22_20_tmp <= r21[20];
r22[20] <= r22_20_tmp;

r22_21_tmp <= r21[21];
r22[21] <= r22_21_tmp;

r22_22_tmp <= r21[22];
r22[22] <= r22_22_tmp;

r22_23_tmp <= r21[23];
r22[23] <= r22_23_tmp;

r22_24_tmp <= r21[24];
r22[24] <= r22_24_tmp;

r22_25_tmp <= r21[25];
r22[25] <= r22_25_tmp;

r22_26_tmp <= r21[26];
r22[26] <= r22_26_tmp;

r22_27_tmp <= r21[27];
r22[27] <= r22_27_tmp;

r22_28_tmp <= r21[28];
r22[28] <= r22_28_tmp;

r22_29_tmp <= r21[29];
r22[29] <= r22_29_tmp;

r22_30_tmp <= r21[30];
r22[30] <= r22_30_tmp;

r22_31_tmp <= r21[31];
r22[31] <= r22_31_tmp;

r22_32_tmp <= r21[32];
r22[32] <= r22_32_tmp;

r22_33_tmp <= r21[33];
r22[33] <= r22_33_tmp;

r22_34_tmp <= r21[34];
r22[34] <= r22_34_tmp;

r22_35_tmp <= r21[35];
r22[35] <= r22_35_tmp;

r22_36_tmp <= r21[36];
r22[36] <= r22_36_tmp;

r22_37_tmp <= r21[37];
r22[37] <= r22_37_tmp;

r22_38_tmp <= r21[38];
r22[38] <= r22_38_tmp;

r22_39_tmp <= r21[39];
r22[39] <= r22_39_tmp;

r22_40_tmp <= r21[40];
r22[40] <= r22_40_tmp;

r22_41_tmp <= r21[41];
r22[41] <= r22_41_tmp;

r22_42_tmp <= r21[42];
r22[42] <= r22_42_tmp;

r22_43_tmp <= r21[43];
r22[43] <= r22_43_tmp;

r22_44_tmp <= r21[44];
r22[44] <= r22_44_tmp;

r22_45_tmp <= r21[45];
r22[45] <= r22_45_tmp;

r22_46_tmp <= r21[46];
r22[46] <= r22_46_tmp;

r22_47_tmp <= r21[47];
r22[47] <= r22_47_tmp;

r22_48_tmp <= r21[48];
r22[48] <= r22_48_tmp;

r22_49_tmp <= r21[49];
r22[49] <= r22_49_tmp;

r22_50_tmp <= r21[50];
r22[50] <= r22_50_tmp;

r22_51_tmp <= r21[51];
r22[51] <= r22_51_tmp;

r22_52_tmp <= r21[52];
r22[52] <= r22_52_tmp;

r22_53_tmp <= r21[53];
r22[53] <= r22_53_tmp;

r22_54_tmp <= r21[54];
r22[54] <= r22_54_tmp;

r22_55_tmp <= r21[55];
r22[55] <= r22_55_tmp;

r22_56_tmp <= r21[56];
r22[56] <= r22_56_tmp;

r22_57_tmp <= r21[57];
r22[57] <= r22_57_tmp;

r22_58_tmp <= r21[58];
r22[58] <= r22_58_tmp;

r22_59_tmp <= r21[59];
r22[59] <= r22_59_tmp;

r22_60_tmp <= r21[60];
r22[60] <= r22_60_tmp;

r22_61_tmp <= r21[61];
r22[61] <= r22_61_tmp;

r22_62_tmp <= r21[62];
r22[62] <= r22_62_tmp;

r22_63_tmp <= r21[63];
r22[63] <= r22_63_tmp;

r22_65_tmp <= r21[65];
r22[65] <= r22_65_tmp;

r22_67_tmp <= r21[67];
r22[67] <= r22_67_tmp;

r22_69_tmp <= r21[69];
r22[69] <= r22_69_tmp;

r22_71_tmp <= r21[71];
r22[71] <= r22_71_tmp;

r22_73_tmp <= r21[73];
r22[73] <= r22_73_tmp;

r22_75_tmp <= r21[75];
r22[75] <= r22_75_tmp;

r22_77_tmp <= r21[77];
r22[77] <= r22_77_tmp;

r22_79_tmp <= r21[79];
r22[79] <= r22_79_tmp;

//--------------------------
//---------layer : 23------------
cmp630_in0 <= r22[9];
cmp630_in1 <= r22[40];
r23[9] <= cmp630_out0;
r23[40] <= cmp630_out1;

cmp631_in0 <= r22[11];
cmp631_in1 <= r22[42];
r23[11] <= cmp631_out0;
r23[42] <= cmp631_out1;

cmp632_in0 <= r22[13];
cmp632_in1 <= r22[44];
r23[13] <= cmp632_out0;
r23[44] <= cmp632_out1;

cmp633_in0 <= r22[15];
cmp633_in1 <= r22[46];
r23[15] <= cmp633_out0;
r23[46] <= cmp633_out1;

cmp634_in0 <= r22[17];
cmp634_in1 <= r22[48];
r23[17] <= cmp634_out0;
r23[48] <= cmp634_out1;

cmp635_in0 <= r22[19];
cmp635_in1 <= r22[50];
r23[19] <= cmp635_out0;
r23[50] <= cmp635_out1;

cmp636_in0 <= r22[21];
cmp636_in1 <= r22[52];
r23[21] <= cmp636_out0;
r23[52] <= cmp636_out1;

cmp637_in0 <= r22[23];
cmp637_in1 <= r22[54];
r23[23] <= cmp637_out0;
r23[54] <= cmp637_out1;

cmp638_in0 <= r22[25];
cmp638_in1 <= r22[56];
r23[25] <= cmp638_out0;
r23[56] <= cmp638_out1;

cmp639_in0 <= r22[27];
cmp639_in1 <= r22[58];
r23[27] <= cmp639_out0;
r23[58] <= cmp639_out1;

cmp640_in0 <= r22[29];
cmp640_in1 <= r22[60];
r23[29] <= cmp640_out0;
r23[60] <= cmp640_out1;

cmp641_in0 <= r22[31];
cmp641_in1 <= r22[62];
r23[31] <= cmp641_out0;
r23[62] <= cmp641_out1;

cmp642_in0 <= r22[33];
cmp642_in1 <= r22[64];
r23[33] <= cmp642_out0;
r23[64] <= cmp642_out1;

cmp643_in0 <= r22[35];
cmp643_in1 <= r22[66];
r23[35] <= cmp643_out0;
r23[66] <= cmp643_out1;

cmp644_in0 <= r22[37];
cmp644_in1 <= r22[68];
r23[37] <= cmp644_out0;
r23[68] <= cmp644_out1;

cmp645_in0 <= r22[39];
cmp645_in1 <= r22[70];
r23[39] <= cmp645_out0;
r23[70] <= cmp645_out1;

r23_0_tmp <= r22[0];
r23[0] <= r23_0_tmp;

r23_1_tmp <= r22[1];
r23[1] <= r23_1_tmp;

r23_2_tmp <= r22[2];
r23[2] <= r23_2_tmp;

r23_3_tmp <= r22[3];
r23[3] <= r23_3_tmp;

r23_4_tmp <= r22[4];
r23[4] <= r23_4_tmp;

r23_5_tmp <= r22[5];
r23[5] <= r23_5_tmp;

r23_6_tmp <= r22[6];
r23[6] <= r23_6_tmp;

r23_7_tmp <= r22[7];
r23[7] <= r23_7_tmp;

r23_8_tmp <= r22[8];
r23[8] <= r23_8_tmp;

r23_10_tmp <= r22[10];
r23[10] <= r23_10_tmp;

r23_12_tmp <= r22[12];
r23[12] <= r23_12_tmp;

r23_14_tmp <= r22[14];
r23[14] <= r23_14_tmp;

r23_16_tmp <= r22[16];
r23[16] <= r23_16_tmp;

r23_18_tmp <= r22[18];
r23[18] <= r23_18_tmp;

r23_20_tmp <= r22[20];
r23[20] <= r23_20_tmp;

r23_22_tmp <= r22[22];
r23[22] <= r23_22_tmp;

r23_24_tmp <= r22[24];
r23[24] <= r23_24_tmp;

r23_26_tmp <= r22[26];
r23[26] <= r23_26_tmp;

r23_28_tmp <= r22[28];
r23[28] <= r23_28_tmp;

r23_30_tmp <= r22[30];
r23[30] <= r23_30_tmp;

r23_32_tmp <= r22[32];
r23[32] <= r23_32_tmp;

r23_34_tmp <= r22[34];
r23[34] <= r23_34_tmp;

r23_36_tmp <= r22[36];
r23[36] <= r23_36_tmp;

r23_38_tmp <= r22[38];
r23[38] <= r23_38_tmp;

r23_41_tmp <= r22[41];
r23[41] <= r23_41_tmp;

r23_43_tmp <= r22[43];
r23[43] <= r23_43_tmp;

r23_45_tmp <= r22[45];
r23[45] <= r23_45_tmp;

r23_47_tmp <= r22[47];
r23[47] <= r23_47_tmp;

r23_49_tmp <= r22[49];
r23[49] <= r23_49_tmp;

r23_51_tmp <= r22[51];
r23[51] <= r23_51_tmp;

r23_53_tmp <= r22[53];
r23[53] <= r23_53_tmp;

r23_55_tmp <= r22[55];
r23[55] <= r23_55_tmp;

r23_57_tmp <= r22[57];
r23[57] <= r23_57_tmp;

r23_59_tmp <= r22[59];
r23[59] <= r23_59_tmp;

r23_61_tmp <= r22[61];
r23[61] <= r23_61_tmp;

r23_63_tmp <= r22[63];
r23[63] <= r23_63_tmp;

r23_65_tmp <= r22[65];
r23[65] <= r23_65_tmp;

r23_67_tmp <= r22[67];
r23[67] <= r23_67_tmp;

r23_69_tmp <= r22[69];
r23[69] <= r23_69_tmp;

r23_71_tmp <= r22[71];
r23[71] <= r23_71_tmp;

r23_72_tmp <= r22[72];
r23[72] <= r23_72_tmp;

r23_73_tmp <= r22[73];
r23[73] <= r23_73_tmp;

r23_74_tmp <= r22[74];
r23[74] <= r23_74_tmp;

r23_75_tmp <= r22[75];
r23[75] <= r23_75_tmp;

r23_76_tmp <= r22[76];
r23[76] <= r23_76_tmp;

r23_77_tmp <= r22[77];
r23[77] <= r23_77_tmp;

r23_78_tmp <= r22[78];
r23[78] <= r23_78_tmp;

r23_79_tmp <= r22[79];
r23[79] <= r23_79_tmp;

r23_80_tmp <= r22[80];
r23[80] <= r23_80_tmp;

//--------------------------
//---------layer : 24------------
cmp646_in0 <= r23[25];
cmp646_in1 <= r23[40];
r24[25] <= cmp646_out0;
r24[40] <= cmp646_out1;

cmp647_in0 <= r23[27];
cmp647_in1 <= r23[42];
r24[27] <= cmp647_out0;
r24[42] <= cmp647_out1;

cmp648_in0 <= r23[29];
cmp648_in1 <= r23[44];
r24[29] <= cmp648_out0;
r24[44] <= cmp648_out1;

cmp649_in0 <= r23[31];
cmp649_in1 <= r23[46];
r24[31] <= cmp649_out0;
r24[46] <= cmp649_out1;

cmp650_in0 <= r23[33];
cmp650_in1 <= r23[48];
r24[33] <= cmp650_out0;
r24[48] <= cmp650_out1;

cmp651_in0 <= r23[35];
cmp651_in1 <= r23[50];
r24[35] <= cmp651_out0;
r24[50] <= cmp651_out1;

cmp652_in0 <= r23[37];
cmp652_in1 <= r23[52];
r24[37] <= cmp652_out0;
r24[52] <= cmp652_out1;

cmp653_in0 <= r23[39];
cmp653_in1 <= r23[54];
r24[39] <= cmp653_out0;
r24[54] <= cmp653_out1;

r24_0_tmp <= r23[0];
r24[0] <= r24_0_tmp;

r24_1_tmp <= r23[1];
r24[1] <= r24_1_tmp;

r24_2_tmp <= r23[2];
r24[2] <= r24_2_tmp;

r24_3_tmp <= r23[3];
r24[3] <= r24_3_tmp;

r24_4_tmp <= r23[4];
r24[4] <= r24_4_tmp;

r24_5_tmp <= r23[5];
r24[5] <= r24_5_tmp;

r24_6_tmp <= r23[6];
r24[6] <= r24_6_tmp;

r24_7_tmp <= r23[7];
r24[7] <= r24_7_tmp;

r24_8_tmp <= r23[8];
r24[8] <= r24_8_tmp;

r24_9_tmp <= r23[9];
r24[9] <= r24_9_tmp;

r24_10_tmp <= r23[10];
r24[10] <= r24_10_tmp;

r24_11_tmp <= r23[11];
r24[11] <= r24_11_tmp;

r24_12_tmp <= r23[12];
r24[12] <= r24_12_tmp;

r24_13_tmp <= r23[13];
r24[13] <= r24_13_tmp;

r24_14_tmp <= r23[14];
r24[14] <= r24_14_tmp;

r24_15_tmp <= r23[15];
r24[15] <= r24_15_tmp;

r24_16_tmp <= r23[16];
r24[16] <= r24_16_tmp;

r24_17_tmp <= r23[17];
r24[17] <= r24_17_tmp;

r24_18_tmp <= r23[18];
r24[18] <= r24_18_tmp;

r24_19_tmp <= r23[19];
r24[19] <= r24_19_tmp;

r24_20_tmp <= r23[20];
r24[20] <= r24_20_tmp;

r24_21_tmp <= r23[21];
r24[21] <= r24_21_tmp;

r24_22_tmp <= r23[22];
r24[22] <= r24_22_tmp;

r24_23_tmp <= r23[23];
r24[23] <= r24_23_tmp;

r24_24_tmp <= r23[24];
r24[24] <= r24_24_tmp;

r24_26_tmp <= r23[26];
r24[26] <= r24_26_tmp;

r24_28_tmp <= r23[28];
r24[28] <= r24_28_tmp;

r24_30_tmp <= r23[30];
r24[30] <= r24_30_tmp;

r24_32_tmp <= r23[32];
r24[32] <= r24_32_tmp;

r24_34_tmp <= r23[34];
r24[34] <= r24_34_tmp;

r24_36_tmp <= r23[36];
r24[36] <= r24_36_tmp;

r24_38_tmp <= r23[38];
r24[38] <= r24_38_tmp;

r24_41_tmp <= r23[41];
r24[41] <= r24_41_tmp;

r24_43_tmp <= r23[43];
r24[43] <= r24_43_tmp;

r24_45_tmp <= r23[45];
r24[45] <= r24_45_tmp;

r24_47_tmp <= r23[47];
r24[47] <= r24_47_tmp;

r24_49_tmp <= r23[49];
r24[49] <= r24_49_tmp;

r24_51_tmp <= r23[51];
r24[51] <= r24_51_tmp;

r24_53_tmp <= r23[53];
r24[53] <= r24_53_tmp;

r24_55_tmp <= r23[55];
r24[55] <= r24_55_tmp;

r24_56_tmp <= r23[56];
r24[56] <= r24_56_tmp;

r24_57_tmp <= r23[57];
r24[57] <= r24_57_tmp;

r24_58_tmp <= r23[58];
r24[58] <= r24_58_tmp;

r24_59_tmp <= r23[59];
r24[59] <= r24_59_tmp;

r24_60_tmp <= r23[60];
r24[60] <= r24_60_tmp;

r24_61_tmp <= r23[61];
r24[61] <= r24_61_tmp;

r24_62_tmp <= r23[62];
r24[62] <= r24_62_tmp;

r24_63_tmp <= r23[63];
r24[63] <= r24_63_tmp;

r24_64_tmp <= r23[64];
r24[64] <= r24_64_tmp;

r24_65_tmp <= r23[65];
r24[65] <= r24_65_tmp;

r24_66_tmp <= r23[66];
r24[66] <= r24_66_tmp;

r24_67_tmp <= r23[67];
r24[67] <= r24_67_tmp;

r24_68_tmp <= r23[68];
r24[68] <= r24_68_tmp;

r24_69_tmp <= r23[69];
r24[69] <= r24_69_tmp;

r24_70_tmp <= r23[70];
r24[70] <= r24_70_tmp;

r24_71_tmp <= r23[71];
r24[71] <= r24_71_tmp;

r24_72_tmp <= r23[72];
r24[72] <= r24_72_tmp;

r24_73_tmp <= r23[73];
r24[73] <= r24_73_tmp;

r24_74_tmp <= r23[74];
r24[74] <= r24_74_tmp;

r24_75_tmp <= r23[75];
r24[75] <= r24_75_tmp;

r24_76_tmp <= r23[76];
r24[76] <= r24_76_tmp;

r24_77_tmp <= r23[77];
r24[77] <= r24_77_tmp;

r24_78_tmp <= r23[78];
r24[78] <= r24_78_tmp;

r24_79_tmp <= r23[79];
r24[79] <= r24_79_tmp;

r24_80_tmp <= r23[80];
r24[80] <= r24_80_tmp;

//--------------------------
//---------layer : 25------------
cmp654_in0 <= r24[33];
cmp654_in1 <= r24[40];
r25[33] <= cmp654_out0;
r25[40] <= cmp654_out1;

cmp655_in0 <= r24[35];
cmp655_in1 <= r24[42];
r25[35] <= cmp655_out0;
r25[42] <= cmp655_out1;

cmp656_in0 <= r24[37];
cmp656_in1 <= r24[44];
r25[37] <= cmp656_out0;
r25[44] <= cmp656_out1;

cmp657_in0 <= r24[39];
cmp657_in1 <= r24[46];
r25[39] <= cmp657_out0;
r25[46] <= cmp657_out1;

r25_0_tmp <= r24[0];
r25[0] <= r25_0_tmp;

r25_1_tmp <= r24[1];
r25[1] <= r25_1_tmp;

r25_2_tmp <= r24[2];
r25[2] <= r25_2_tmp;

r25_3_tmp <= r24[3];
r25[3] <= r25_3_tmp;

r25_4_tmp <= r24[4];
r25[4] <= r25_4_tmp;

r25_5_tmp <= r24[5];
r25[5] <= r25_5_tmp;

r25_6_tmp <= r24[6];
r25[6] <= r25_6_tmp;

r25_7_tmp <= r24[7];
r25[7] <= r25_7_tmp;

r25_8_tmp <= r24[8];
r25[8] <= r25_8_tmp;

r25_9_tmp <= r24[9];
r25[9] <= r25_9_tmp;

r25_10_tmp <= r24[10];
r25[10] <= r25_10_tmp;

r25_11_tmp <= r24[11];
r25[11] <= r25_11_tmp;

r25_12_tmp <= r24[12];
r25[12] <= r25_12_tmp;

r25_13_tmp <= r24[13];
r25[13] <= r25_13_tmp;

r25_14_tmp <= r24[14];
r25[14] <= r25_14_tmp;

r25_15_tmp <= r24[15];
r25[15] <= r25_15_tmp;

r25_16_tmp <= r24[16];
r25[16] <= r25_16_tmp;

r25_17_tmp <= r24[17];
r25[17] <= r25_17_tmp;

r25_18_tmp <= r24[18];
r25[18] <= r25_18_tmp;

r25_19_tmp <= r24[19];
r25[19] <= r25_19_tmp;

r25_20_tmp <= r24[20];
r25[20] <= r25_20_tmp;

r25_21_tmp <= r24[21];
r25[21] <= r25_21_tmp;

r25_22_tmp <= r24[22];
r25[22] <= r25_22_tmp;

r25_23_tmp <= r24[23];
r25[23] <= r25_23_tmp;

r25_24_tmp <= r24[24];
r25[24] <= r25_24_tmp;

r25_25_tmp <= r24[25];
r25[25] <= r25_25_tmp;

r25_26_tmp <= r24[26];
r25[26] <= r25_26_tmp;

r25_27_tmp <= r24[27];
r25[27] <= r25_27_tmp;

r25_28_tmp <= r24[28];
r25[28] <= r25_28_tmp;

r25_29_tmp <= r24[29];
r25[29] <= r25_29_tmp;

r25_30_tmp <= r24[30];
r25[30] <= r25_30_tmp;

r25_31_tmp <= r24[31];
r25[31] <= r25_31_tmp;

r25_32_tmp <= r24[32];
r25[32] <= r25_32_tmp;

r25_34_tmp <= r24[34];
r25[34] <= r25_34_tmp;

r25_36_tmp <= r24[36];
r25[36] <= r25_36_tmp;

r25_38_tmp <= r24[38];
r25[38] <= r25_38_tmp;

r25_41_tmp <= r24[41];
r25[41] <= r25_41_tmp;

r25_43_tmp <= r24[43];
r25[43] <= r25_43_tmp;

r25_45_tmp <= r24[45];
r25[45] <= r25_45_tmp;

r25_47_tmp <= r24[47];
r25[47] <= r25_47_tmp;

r25_48_tmp <= r24[48];
r25[48] <= r25_48_tmp;

r25_49_tmp <= r24[49];
r25[49] <= r25_49_tmp;

r25_50_tmp <= r24[50];
r25[50] <= r25_50_tmp;

r25_51_tmp <= r24[51];
r25[51] <= r25_51_tmp;

r25_52_tmp <= r24[52];
r25[52] <= r25_52_tmp;

r25_53_tmp <= r24[53];
r25[53] <= r25_53_tmp;

r25_54_tmp <= r24[54];
r25[54] <= r25_54_tmp;

r25_55_tmp <= r24[55];
r25[55] <= r25_55_tmp;

r25_56_tmp <= r24[56];
r25[56] <= r25_56_tmp;

r25_57_tmp <= r24[57];
r25[57] <= r25_57_tmp;

r25_58_tmp <= r24[58];
r25[58] <= r25_58_tmp;

r25_59_tmp <= r24[59];
r25[59] <= r25_59_tmp;

r25_60_tmp <= r24[60];
r25[60] <= r25_60_tmp;

r25_61_tmp <= r24[61];
r25[61] <= r25_61_tmp;

r25_62_tmp <= r24[62];
r25[62] <= r25_62_tmp;

r25_63_tmp <= r24[63];
r25[63] <= r25_63_tmp;

r25_64_tmp <= r24[64];
r25[64] <= r25_64_tmp;

r25_65_tmp <= r24[65];
r25[65] <= r25_65_tmp;

r25_66_tmp <= r24[66];
r25[66] <= r25_66_tmp;

r25_67_tmp <= r24[67];
r25[67] <= r25_67_tmp;

r25_68_tmp <= r24[68];
r25[68] <= r25_68_tmp;

r25_69_tmp <= r24[69];
r25[69] <= r25_69_tmp;

r25_70_tmp <= r24[70];
r25[70] <= r25_70_tmp;

r25_71_tmp <= r24[71];
r25[71] <= r25_71_tmp;

r25_72_tmp <= r24[72];
r25[72] <= r25_72_tmp;

r25_73_tmp <= r24[73];
r25[73] <= r25_73_tmp;

r25_74_tmp <= r24[74];
r25[74] <= r25_74_tmp;

r25_75_tmp <= r24[75];
r25[75] <= r25_75_tmp;

r25_76_tmp <= r24[76];
r25[76] <= r25_76_tmp;

r25_77_tmp <= r24[77];
r25[77] <= r25_77_tmp;

r25_78_tmp <= r24[78];
r25[78] <= r25_78_tmp;

r25_79_tmp <= r24[79];
r25[79] <= r25_79_tmp;

r25_80_tmp <= r24[80];
r25[80] <= r25_80_tmp;

//--------------------------
//---------layer : 26------------
cmp658_in0 <= r25[37];
cmp658_in1 <= r25[40];
r26[37] <= cmp658_out0;
r26[40] <= cmp658_out1;

cmp659_in0 <= r25[39];
cmp659_in1 <= r25[42];
r26[39] <= cmp659_out0;
r26[42] <= cmp659_out1;

r26_0_tmp <= r25[0];
r26[0] <= r26_0_tmp;

r26_1_tmp <= r25[1];
r26[1] <= r26_1_tmp;

r26_2_tmp <= r25[2];
r26[2] <= r26_2_tmp;

r26_3_tmp <= r25[3];
r26[3] <= r26_3_tmp;

r26_4_tmp <= r25[4];
r26[4] <= r26_4_tmp;

r26_5_tmp <= r25[5];
r26[5] <= r26_5_tmp;

r26_6_tmp <= r25[6];
r26[6] <= r26_6_tmp;

r26_7_tmp <= r25[7];
r26[7] <= r26_7_tmp;

r26_8_tmp <= r25[8];
r26[8] <= r26_8_tmp;

r26_9_tmp <= r25[9];
r26[9] <= r26_9_tmp;

r26_10_tmp <= r25[10];
r26[10] <= r26_10_tmp;

r26_11_tmp <= r25[11];
r26[11] <= r26_11_tmp;

r26_12_tmp <= r25[12];
r26[12] <= r26_12_tmp;

r26_13_tmp <= r25[13];
r26[13] <= r26_13_tmp;

r26_14_tmp <= r25[14];
r26[14] <= r26_14_tmp;

r26_15_tmp <= r25[15];
r26[15] <= r26_15_tmp;

r26_16_tmp <= r25[16];
r26[16] <= r26_16_tmp;

r26_17_tmp <= r25[17];
r26[17] <= r26_17_tmp;

r26_18_tmp <= r25[18];
r26[18] <= r26_18_tmp;

r26_19_tmp <= r25[19];
r26[19] <= r26_19_tmp;

r26_20_tmp <= r25[20];
r26[20] <= r26_20_tmp;

r26_21_tmp <= r25[21];
r26[21] <= r26_21_tmp;

r26_22_tmp <= r25[22];
r26[22] <= r26_22_tmp;

r26_23_tmp <= r25[23];
r26[23] <= r26_23_tmp;

r26_24_tmp <= r25[24];
r26[24] <= r26_24_tmp;

r26_25_tmp <= r25[25];
r26[25] <= r26_25_tmp;

r26_26_tmp <= r25[26];
r26[26] <= r26_26_tmp;

r26_27_tmp <= r25[27];
r26[27] <= r26_27_tmp;

r26_28_tmp <= r25[28];
r26[28] <= r26_28_tmp;

r26_29_tmp <= r25[29];
r26[29] <= r26_29_tmp;

r26_30_tmp <= r25[30];
r26[30] <= r26_30_tmp;

r26_31_tmp <= r25[31];
r26[31] <= r26_31_tmp;

r26_32_tmp <= r25[32];
r26[32] <= r26_32_tmp;

r26_33_tmp <= r25[33];
r26[33] <= r26_33_tmp;

r26_34_tmp <= r25[34];
r26[34] <= r26_34_tmp;

r26_35_tmp <= r25[35];
r26[35] <= r26_35_tmp;

r26_36_tmp <= r25[36];
r26[36] <= r26_36_tmp;

r26_38_tmp <= r25[38];
r26[38] <= r26_38_tmp;

r26_41_tmp <= r25[41];
r26[41] <= r26_41_tmp;

r26_43_tmp <= r25[43];
r26[43] <= r26_43_tmp;

r26_44_tmp <= r25[44];
r26[44] <= r26_44_tmp;

r26_45_tmp <= r25[45];
r26[45] <= r26_45_tmp;

r26_46_tmp <= r25[46];
r26[46] <= r26_46_tmp;

r26_47_tmp <= r25[47];
r26[47] <= r26_47_tmp;

r26_48_tmp <= r25[48];
r26[48] <= r26_48_tmp;

r26_49_tmp <= r25[49];
r26[49] <= r26_49_tmp;

r26_50_tmp <= r25[50];
r26[50] <= r26_50_tmp;

r26_51_tmp <= r25[51];
r26[51] <= r26_51_tmp;

r26_52_tmp <= r25[52];
r26[52] <= r26_52_tmp;

r26_53_tmp <= r25[53];
r26[53] <= r26_53_tmp;

r26_54_tmp <= r25[54];
r26[54] <= r26_54_tmp;

r26_55_tmp <= r25[55];
r26[55] <= r26_55_tmp;

r26_56_tmp <= r25[56];
r26[56] <= r26_56_tmp;

r26_57_tmp <= r25[57];
r26[57] <= r26_57_tmp;

r26_58_tmp <= r25[58];
r26[58] <= r26_58_tmp;

r26_59_tmp <= r25[59];
r26[59] <= r26_59_tmp;

r26_60_tmp <= r25[60];
r26[60] <= r26_60_tmp;

r26_61_tmp <= r25[61];
r26[61] <= r26_61_tmp;

r26_62_tmp <= r25[62];
r26[62] <= r26_62_tmp;

r26_63_tmp <= r25[63];
r26[63] <= r26_63_tmp;

r26_64_tmp <= r25[64];
r26[64] <= r26_64_tmp;

r26_65_tmp <= r25[65];
r26[65] <= r26_65_tmp;

r26_66_tmp <= r25[66];
r26[66] <= r26_66_tmp;

r26_67_tmp <= r25[67];
r26[67] <= r26_67_tmp;

r26_68_tmp <= r25[68];
r26[68] <= r26_68_tmp;

r26_69_tmp <= r25[69];
r26[69] <= r26_69_tmp;

r26_70_tmp <= r25[70];
r26[70] <= r26_70_tmp;

r26_71_tmp <= r25[71];
r26[71] <= r26_71_tmp;

r26_72_tmp <= r25[72];
r26[72] <= r26_72_tmp;

r26_73_tmp <= r25[73];
r26[73] <= r26_73_tmp;

r26_74_tmp <= r25[74];
r26[74] <= r26_74_tmp;

r26_75_tmp <= r25[75];
r26[75] <= r26_75_tmp;

r26_76_tmp <= r25[76];
r26[76] <= r26_76_tmp;

r26_77_tmp <= r25[77];
r26[77] <= r26_77_tmp;

r26_78_tmp <= r25[78];
r26[78] <= r26_78_tmp;

r26_79_tmp <= r25[79];
r26[79] <= r26_79_tmp;

r26_80_tmp <= r25[80];
r26[80] <= r26_80_tmp;

//--------------------------
//---------layer : 27------------
cmp660_in0 <= r26[39];
cmp660_in1 <= r26[40];
r27[39] <= cmp660_out0;
r27[40] <= cmp660_out1;

r27_0_tmp <= r26[0];
r27[0] <= r27_0_tmp;

r27_1_tmp <= r26[1];
r27[1] <= r27_1_tmp;

r27_2_tmp <= r26[2];
r27[2] <= r27_2_tmp;

r27_3_tmp <= r26[3];
r27[3] <= r27_3_tmp;

r27_4_tmp <= r26[4];
r27[4] <= r27_4_tmp;

r27_5_tmp <= r26[5];
r27[5] <= r27_5_tmp;

r27_6_tmp <= r26[6];
r27[6] <= r27_6_tmp;

r27_7_tmp <= r26[7];
r27[7] <= r27_7_tmp;

r27_8_tmp <= r26[8];
r27[8] <= r27_8_tmp;

r27_9_tmp <= r26[9];
r27[9] <= r27_9_tmp;

r27_10_tmp <= r26[10];
r27[10] <= r27_10_tmp;

r27_11_tmp <= r26[11];
r27[11] <= r27_11_tmp;

r27_12_tmp <= r26[12];
r27[12] <= r27_12_tmp;

r27_13_tmp <= r26[13];
r27[13] <= r27_13_tmp;

r27_14_tmp <= r26[14];
r27[14] <= r27_14_tmp;

r27_15_tmp <= r26[15];
r27[15] <= r27_15_tmp;

r27_16_tmp <= r26[16];
r27[16] <= r27_16_tmp;

r27_17_tmp <= r26[17];
r27[17] <= r27_17_tmp;

r27_18_tmp <= r26[18];
r27[18] <= r27_18_tmp;

r27_19_tmp <= r26[19];
r27[19] <= r27_19_tmp;

r27_20_tmp <= r26[20];
r27[20] <= r27_20_tmp;

r27_21_tmp <= r26[21];
r27[21] <= r27_21_tmp;

r27_22_tmp <= r26[22];
r27[22] <= r27_22_tmp;

r27_23_tmp <= r26[23];
r27[23] <= r27_23_tmp;

r27_24_tmp <= r26[24];
r27[24] <= r27_24_tmp;

r27_25_tmp <= r26[25];
r27[25] <= r27_25_tmp;

r27_26_tmp <= r26[26];
r27[26] <= r27_26_tmp;

r27_27_tmp <= r26[27];
r27[27] <= r27_27_tmp;

r27_28_tmp <= r26[28];
r27[28] <= r27_28_tmp;

r27_29_tmp <= r26[29];
r27[29] <= r27_29_tmp;

r27_30_tmp <= r26[30];
r27[30] <= r27_30_tmp;

r27_31_tmp <= r26[31];
r27[31] <= r27_31_tmp;

r27_32_tmp <= r26[32];
r27[32] <= r27_32_tmp;

r27_33_tmp <= r26[33];
r27[33] <= r27_33_tmp;

r27_34_tmp <= r26[34];
r27[34] <= r27_34_tmp;

r27_35_tmp <= r26[35];
r27[35] <= r27_35_tmp;

r27_36_tmp <= r26[36];
r27[36] <= r27_36_tmp;

r27_37_tmp <= r26[37];
r27[37] <= r27_37_tmp;

r27_38_tmp <= r26[38];
r27[38] <= r27_38_tmp;

r27_41_tmp <= r26[41];
r27[41] <= r27_41_tmp;

r27_42_tmp <= r26[42];
r27[42] <= r27_42_tmp;

r27_43_tmp <= r26[43];
r27[43] <= r27_43_tmp;

r27_44_tmp <= r26[44];
r27[44] <= r27_44_tmp;

r27_45_tmp <= r26[45];
r27[45] <= r27_45_tmp;

r27_46_tmp <= r26[46];
r27[46] <= r27_46_tmp;

r27_47_tmp <= r26[47];
r27[47] <= r27_47_tmp;

r27_48_tmp <= r26[48];
r27[48] <= r27_48_tmp;

r27_49_tmp <= r26[49];
r27[49] <= r27_49_tmp;

r27_50_tmp <= r26[50];
r27[50] <= r27_50_tmp;

r27_51_tmp <= r26[51];
r27[51] <= r27_51_tmp;

r27_52_tmp <= r26[52];
r27[52] <= r27_52_tmp;

r27_53_tmp <= r26[53];
r27[53] <= r27_53_tmp;

r27_54_tmp <= r26[54];
r27[54] <= r27_54_tmp;

r27_55_tmp <= r26[55];
r27[55] <= r27_55_tmp;

r27_56_tmp <= r26[56];
r27[56] <= r27_56_tmp;

r27_57_tmp <= r26[57];
r27[57] <= r27_57_tmp;

r27_58_tmp <= r26[58];
r27[58] <= r27_58_tmp;

r27_59_tmp <= r26[59];
r27[59] <= r27_59_tmp;

r27_60_tmp <= r26[60];
r27[60] <= r27_60_tmp;

r27_61_tmp <= r26[61];
r27[61] <= r27_61_tmp;

r27_62_tmp <= r26[62];
r27[62] <= r27_62_tmp;

r27_63_tmp <= r26[63];
r27[63] <= r27_63_tmp;

r27_64_tmp <= r26[64];
r27[64] <= r27_64_tmp;

r27_65_tmp <= r26[65];
r27[65] <= r27_65_tmp;

r27_66_tmp <= r26[66];
r27[66] <= r27_66_tmp;

r27_67_tmp <= r26[67];
r27[67] <= r27_67_tmp;

r27_68_tmp <= r26[68];
r27[68] <= r27_68_tmp;

r27_69_tmp <= r26[69];
r27[69] <= r27_69_tmp;

r27_70_tmp <= r26[70];
r27[70] <= r27_70_tmp;

r27_71_tmp <= r26[71];
r27[71] <= r27_71_tmp;

r27_72_tmp <= r26[72];
r27[72] <= r27_72_tmp;

r27_73_tmp <= r26[73];
r27[73] <= r27_73_tmp;

r27_74_tmp <= r26[74];
r27[74] <= r27_74_tmp;

r27_75_tmp <= r26[75];
r27[75] <= r27_75_tmp;

r27_76_tmp <= r26[76];
r27[76] <= r27_76_tmp;

r27_77_tmp <= r26[77];
r27[77] <= r27_77_tmp;

r27_78_tmp <= r26[78];
r27[78] <= r27_78_tmp;

r27_79_tmp <= r26[79];
r27[79] <= r27_79_tmp;

r27_80_tmp <= r26[80];
r27[80] <= r27_80_tmp;

//--------------------------
end
//-------------------Comparator module connect-------------------------------
cmp cmp0 (.in0(cmp0_in0), .in1(cmp0_in1), .out0(cmp0_out0), .out1(cmp0_out1));
cmp cmp1 (.in0(cmp1_in0), .in1(cmp1_in1), .out0(cmp1_out0), .out1(cmp1_out1));
cmp cmp2 (.in0(cmp2_in0), .in1(cmp2_in1), .out0(cmp2_out0), .out1(cmp2_out1));
cmp cmp3 (.in0(cmp3_in0), .in1(cmp3_in1), .out0(cmp3_out0), .out1(cmp3_out1));
cmp cmp4 (.in0(cmp4_in0), .in1(cmp4_in1), .out0(cmp4_out0), .out1(cmp4_out1));
cmp cmp5 (.in0(cmp5_in0), .in1(cmp5_in1), .out0(cmp5_out0), .out1(cmp5_out1));
cmp cmp6 (.in0(cmp6_in0), .in1(cmp6_in1), .out0(cmp6_out0), .out1(cmp6_out1));
cmp cmp7 (.in0(cmp7_in0), .in1(cmp7_in1), .out0(cmp7_out0), .out1(cmp7_out1));
cmp cmp8 (.in0(cmp8_in0), .in1(cmp8_in1), .out0(cmp8_out0), .out1(cmp8_out1));
cmp cmp9 (.in0(cmp9_in0), .in1(cmp9_in1), .out0(cmp9_out0), .out1(cmp9_out1));
cmp cmp10 (.in0(cmp10_in0), .in1(cmp10_in1), .out0(cmp10_out0), .out1(cmp10_out1));
cmp cmp11 (.in0(cmp11_in0), .in1(cmp11_in1), .out0(cmp11_out0), .out1(cmp11_out1));
cmp cmp12 (.in0(cmp12_in0), .in1(cmp12_in1), .out0(cmp12_out0), .out1(cmp12_out1));
cmp cmp13 (.in0(cmp13_in0), .in1(cmp13_in1), .out0(cmp13_out0), .out1(cmp13_out1));
cmp cmp14 (.in0(cmp14_in0), .in1(cmp14_in1), .out0(cmp14_out0), .out1(cmp14_out1));
cmp cmp15 (.in0(cmp15_in0), .in1(cmp15_in1), .out0(cmp15_out0), .out1(cmp15_out1));
cmp cmp16 (.in0(cmp16_in0), .in1(cmp16_in1), .out0(cmp16_out0), .out1(cmp16_out1));
cmp cmp17 (.in0(cmp17_in0), .in1(cmp17_in1), .out0(cmp17_out0), .out1(cmp17_out1));
cmp cmp18 (.in0(cmp18_in0), .in1(cmp18_in1), .out0(cmp18_out0), .out1(cmp18_out1));
cmp cmp19 (.in0(cmp19_in0), .in1(cmp19_in1), .out0(cmp19_out0), .out1(cmp19_out1));
cmp cmp20 (.in0(cmp20_in0), .in1(cmp20_in1), .out0(cmp20_out0), .out1(cmp20_out1));
cmp cmp21 (.in0(cmp21_in0), .in1(cmp21_in1), .out0(cmp21_out0), .out1(cmp21_out1));
cmp cmp22 (.in0(cmp22_in0), .in1(cmp22_in1), .out0(cmp22_out0), .out1(cmp22_out1));
cmp cmp23 (.in0(cmp23_in0), .in1(cmp23_in1), .out0(cmp23_out0), .out1(cmp23_out1));
cmp cmp24 (.in0(cmp24_in0), .in1(cmp24_in1), .out0(cmp24_out0), .out1(cmp24_out1));
cmp cmp25 (.in0(cmp25_in0), .in1(cmp25_in1), .out0(cmp25_out0), .out1(cmp25_out1));
cmp cmp26 (.in0(cmp26_in0), .in1(cmp26_in1), .out0(cmp26_out0), .out1(cmp26_out1));
cmp cmp27 (.in0(cmp27_in0), .in1(cmp27_in1), .out0(cmp27_out0), .out1(cmp27_out1));
cmp cmp28 (.in0(cmp28_in0), .in1(cmp28_in1), .out0(cmp28_out0), .out1(cmp28_out1));
cmp cmp29 (.in0(cmp29_in0), .in1(cmp29_in1), .out0(cmp29_out0), .out1(cmp29_out1));
cmp cmp30 (.in0(cmp30_in0), .in1(cmp30_in1), .out0(cmp30_out0), .out1(cmp30_out1));
cmp cmp31 (.in0(cmp31_in0), .in1(cmp31_in1), .out0(cmp31_out0), .out1(cmp31_out1));
cmp cmp32 (.in0(cmp32_in0), .in1(cmp32_in1), .out0(cmp32_out0), .out1(cmp32_out1));
cmp cmp33 (.in0(cmp33_in0), .in1(cmp33_in1), .out0(cmp33_out0), .out1(cmp33_out1));
cmp cmp34 (.in0(cmp34_in0), .in1(cmp34_in1), .out0(cmp34_out0), .out1(cmp34_out1));
cmp cmp35 (.in0(cmp35_in0), .in1(cmp35_in1), .out0(cmp35_out0), .out1(cmp35_out1));
cmp cmp36 (.in0(cmp36_in0), .in1(cmp36_in1), .out0(cmp36_out0), .out1(cmp36_out1));
cmp cmp37 (.in0(cmp37_in0), .in1(cmp37_in1), .out0(cmp37_out0), .out1(cmp37_out1));
cmp cmp38 (.in0(cmp38_in0), .in1(cmp38_in1), .out0(cmp38_out0), .out1(cmp38_out1));
cmp cmp39 (.in0(cmp39_in0), .in1(cmp39_in1), .out0(cmp39_out0), .out1(cmp39_out1));
cmp cmp40 (.in0(cmp40_in0), .in1(cmp40_in1), .out0(cmp40_out0), .out1(cmp40_out1));
cmp cmp41 (.in0(cmp41_in0), .in1(cmp41_in1), .out0(cmp41_out0), .out1(cmp41_out1));
cmp cmp42 (.in0(cmp42_in0), .in1(cmp42_in1), .out0(cmp42_out0), .out1(cmp42_out1));
cmp cmp43 (.in0(cmp43_in0), .in1(cmp43_in1), .out0(cmp43_out0), .out1(cmp43_out1));
cmp cmp44 (.in0(cmp44_in0), .in1(cmp44_in1), .out0(cmp44_out0), .out1(cmp44_out1));
cmp cmp45 (.in0(cmp45_in0), .in1(cmp45_in1), .out0(cmp45_out0), .out1(cmp45_out1));
cmp cmp46 (.in0(cmp46_in0), .in1(cmp46_in1), .out0(cmp46_out0), .out1(cmp46_out1));
cmp cmp47 (.in0(cmp47_in0), .in1(cmp47_in1), .out0(cmp47_out0), .out1(cmp47_out1));
cmp cmp48 (.in0(cmp48_in0), .in1(cmp48_in1), .out0(cmp48_out0), .out1(cmp48_out1));
cmp cmp49 (.in0(cmp49_in0), .in1(cmp49_in1), .out0(cmp49_out0), .out1(cmp49_out1));
cmp cmp50 (.in0(cmp50_in0), .in1(cmp50_in1), .out0(cmp50_out0), .out1(cmp50_out1));
cmp cmp51 (.in0(cmp51_in0), .in1(cmp51_in1), .out0(cmp51_out0), .out1(cmp51_out1));
cmp cmp52 (.in0(cmp52_in0), .in1(cmp52_in1), .out0(cmp52_out0), .out1(cmp52_out1));
cmp cmp53 (.in0(cmp53_in0), .in1(cmp53_in1), .out0(cmp53_out0), .out1(cmp53_out1));
cmp cmp54 (.in0(cmp54_in0), .in1(cmp54_in1), .out0(cmp54_out0), .out1(cmp54_out1));
cmp cmp55 (.in0(cmp55_in0), .in1(cmp55_in1), .out0(cmp55_out0), .out1(cmp55_out1));
cmp cmp56 (.in0(cmp56_in0), .in1(cmp56_in1), .out0(cmp56_out0), .out1(cmp56_out1));
cmp cmp57 (.in0(cmp57_in0), .in1(cmp57_in1), .out0(cmp57_out0), .out1(cmp57_out1));
cmp cmp58 (.in0(cmp58_in0), .in1(cmp58_in1), .out0(cmp58_out0), .out1(cmp58_out1));
cmp cmp59 (.in0(cmp59_in0), .in1(cmp59_in1), .out0(cmp59_out0), .out1(cmp59_out1));
cmp cmp60 (.in0(cmp60_in0), .in1(cmp60_in1), .out0(cmp60_out0), .out1(cmp60_out1));
cmp cmp61 (.in0(cmp61_in0), .in1(cmp61_in1), .out0(cmp61_out0), .out1(cmp61_out1));
cmp cmp62 (.in0(cmp62_in0), .in1(cmp62_in1), .out0(cmp62_out0), .out1(cmp62_out1));
cmp cmp63 (.in0(cmp63_in0), .in1(cmp63_in1), .out0(cmp63_out0), .out1(cmp63_out1));
cmp cmp64 (.in0(cmp64_in0), .in1(cmp64_in1), .out0(cmp64_out0), .out1(cmp64_out1));
cmp cmp65 (.in0(cmp65_in0), .in1(cmp65_in1), .out0(cmp65_out0), .out1(cmp65_out1));
cmp cmp66 (.in0(cmp66_in0), .in1(cmp66_in1), .out0(cmp66_out0), .out1(cmp66_out1));
cmp cmp67 (.in0(cmp67_in0), .in1(cmp67_in1), .out0(cmp67_out0), .out1(cmp67_out1));
cmp cmp68 (.in0(cmp68_in0), .in1(cmp68_in1), .out0(cmp68_out0), .out1(cmp68_out1));
cmp cmp69 (.in0(cmp69_in0), .in1(cmp69_in1), .out0(cmp69_out0), .out1(cmp69_out1));
cmp cmp70 (.in0(cmp70_in0), .in1(cmp70_in1), .out0(cmp70_out0), .out1(cmp70_out1));
cmp cmp71 (.in0(cmp71_in0), .in1(cmp71_in1), .out0(cmp71_out0), .out1(cmp71_out1));
cmp cmp72 (.in0(cmp72_in0), .in1(cmp72_in1), .out0(cmp72_out0), .out1(cmp72_out1));
cmp cmp73 (.in0(cmp73_in0), .in1(cmp73_in1), .out0(cmp73_out0), .out1(cmp73_out1));
cmp cmp74 (.in0(cmp74_in0), .in1(cmp74_in1), .out0(cmp74_out0), .out1(cmp74_out1));
cmp cmp75 (.in0(cmp75_in0), .in1(cmp75_in1), .out0(cmp75_out0), .out1(cmp75_out1));
cmp cmp76 (.in0(cmp76_in0), .in1(cmp76_in1), .out0(cmp76_out0), .out1(cmp76_out1));
cmp cmp77 (.in0(cmp77_in0), .in1(cmp77_in1), .out0(cmp77_out0), .out1(cmp77_out1));
cmp cmp78 (.in0(cmp78_in0), .in1(cmp78_in1), .out0(cmp78_out0), .out1(cmp78_out1));
cmp cmp79 (.in0(cmp79_in0), .in1(cmp79_in1), .out0(cmp79_out0), .out1(cmp79_out1));
cmp cmp80 (.in0(cmp80_in0), .in1(cmp80_in1), .out0(cmp80_out0), .out1(cmp80_out1));
cmp cmp81 (.in0(cmp81_in0), .in1(cmp81_in1), .out0(cmp81_out0), .out1(cmp81_out1));
cmp cmp82 (.in0(cmp82_in0), .in1(cmp82_in1), .out0(cmp82_out0), .out1(cmp82_out1));
cmp cmp83 (.in0(cmp83_in0), .in1(cmp83_in1), .out0(cmp83_out0), .out1(cmp83_out1));
cmp cmp84 (.in0(cmp84_in0), .in1(cmp84_in1), .out0(cmp84_out0), .out1(cmp84_out1));
cmp cmp85 (.in0(cmp85_in0), .in1(cmp85_in1), .out0(cmp85_out0), .out1(cmp85_out1));
cmp cmp86 (.in0(cmp86_in0), .in1(cmp86_in1), .out0(cmp86_out0), .out1(cmp86_out1));
cmp cmp87 (.in0(cmp87_in0), .in1(cmp87_in1), .out0(cmp87_out0), .out1(cmp87_out1));
cmp cmp88 (.in0(cmp88_in0), .in1(cmp88_in1), .out0(cmp88_out0), .out1(cmp88_out1));
cmp cmp89 (.in0(cmp89_in0), .in1(cmp89_in1), .out0(cmp89_out0), .out1(cmp89_out1));
cmp cmp90 (.in0(cmp90_in0), .in1(cmp90_in1), .out0(cmp90_out0), .out1(cmp90_out1));
cmp cmp91 (.in0(cmp91_in0), .in1(cmp91_in1), .out0(cmp91_out0), .out1(cmp91_out1));
cmp cmp92 (.in0(cmp92_in0), .in1(cmp92_in1), .out0(cmp92_out0), .out1(cmp92_out1));
cmp cmp93 (.in0(cmp93_in0), .in1(cmp93_in1), .out0(cmp93_out0), .out1(cmp93_out1));
cmp cmp94 (.in0(cmp94_in0), .in1(cmp94_in1), .out0(cmp94_out0), .out1(cmp94_out1));
cmp cmp95 (.in0(cmp95_in0), .in1(cmp95_in1), .out0(cmp95_out0), .out1(cmp95_out1));
cmp cmp96 (.in0(cmp96_in0), .in1(cmp96_in1), .out0(cmp96_out0), .out1(cmp96_out1));
cmp cmp97 (.in0(cmp97_in0), .in1(cmp97_in1), .out0(cmp97_out0), .out1(cmp97_out1));
cmp cmp98 (.in0(cmp98_in0), .in1(cmp98_in1), .out0(cmp98_out0), .out1(cmp98_out1));
cmp cmp99 (.in0(cmp99_in0), .in1(cmp99_in1), .out0(cmp99_out0), .out1(cmp99_out1));
cmp cmp100 (.in0(cmp100_in0), .in1(cmp100_in1), .out0(cmp100_out0), .out1(cmp100_out1));
cmp cmp101 (.in0(cmp101_in0), .in1(cmp101_in1), .out0(cmp101_out0), .out1(cmp101_out1));
cmp cmp102 (.in0(cmp102_in0), .in1(cmp102_in1), .out0(cmp102_out0), .out1(cmp102_out1));
cmp cmp103 (.in0(cmp103_in0), .in1(cmp103_in1), .out0(cmp103_out0), .out1(cmp103_out1));
cmp cmp104 (.in0(cmp104_in0), .in1(cmp104_in1), .out0(cmp104_out0), .out1(cmp104_out1));
cmp cmp105 (.in0(cmp105_in0), .in1(cmp105_in1), .out0(cmp105_out0), .out1(cmp105_out1));
cmp cmp106 (.in0(cmp106_in0), .in1(cmp106_in1), .out0(cmp106_out0), .out1(cmp106_out1));
cmp cmp107 (.in0(cmp107_in0), .in1(cmp107_in1), .out0(cmp107_out0), .out1(cmp107_out1));
cmp cmp108 (.in0(cmp108_in0), .in1(cmp108_in1), .out0(cmp108_out0), .out1(cmp108_out1));
cmp cmp109 (.in0(cmp109_in0), .in1(cmp109_in1), .out0(cmp109_out0), .out1(cmp109_out1));
cmp cmp110 (.in0(cmp110_in0), .in1(cmp110_in1), .out0(cmp110_out0), .out1(cmp110_out1));
cmp cmp111 (.in0(cmp111_in0), .in1(cmp111_in1), .out0(cmp111_out0), .out1(cmp111_out1));
cmp cmp112 (.in0(cmp112_in0), .in1(cmp112_in1), .out0(cmp112_out0), .out1(cmp112_out1));
cmp cmp113 (.in0(cmp113_in0), .in1(cmp113_in1), .out0(cmp113_out0), .out1(cmp113_out1));
cmp cmp114 (.in0(cmp114_in0), .in1(cmp114_in1), .out0(cmp114_out0), .out1(cmp114_out1));
cmp cmp115 (.in0(cmp115_in0), .in1(cmp115_in1), .out0(cmp115_out0), .out1(cmp115_out1));
cmp cmp116 (.in0(cmp116_in0), .in1(cmp116_in1), .out0(cmp116_out0), .out1(cmp116_out1));
cmp cmp117 (.in0(cmp117_in0), .in1(cmp117_in1), .out0(cmp117_out0), .out1(cmp117_out1));
cmp cmp118 (.in0(cmp118_in0), .in1(cmp118_in1), .out0(cmp118_out0), .out1(cmp118_out1));
cmp cmp119 (.in0(cmp119_in0), .in1(cmp119_in1), .out0(cmp119_out0), .out1(cmp119_out1));
cmp cmp120 (.in0(cmp120_in0), .in1(cmp120_in1), .out0(cmp120_out0), .out1(cmp120_out1));
cmp cmp121 (.in0(cmp121_in0), .in1(cmp121_in1), .out0(cmp121_out0), .out1(cmp121_out1));
cmp cmp122 (.in0(cmp122_in0), .in1(cmp122_in1), .out0(cmp122_out0), .out1(cmp122_out1));
cmp cmp123 (.in0(cmp123_in0), .in1(cmp123_in1), .out0(cmp123_out0), .out1(cmp123_out1));
cmp cmp124 (.in0(cmp124_in0), .in1(cmp124_in1), .out0(cmp124_out0), .out1(cmp124_out1));
cmp cmp125 (.in0(cmp125_in0), .in1(cmp125_in1), .out0(cmp125_out0), .out1(cmp125_out1));
cmp cmp126 (.in0(cmp126_in0), .in1(cmp126_in1), .out0(cmp126_out0), .out1(cmp126_out1));
cmp cmp127 (.in0(cmp127_in0), .in1(cmp127_in1), .out0(cmp127_out0), .out1(cmp127_out1));
cmp cmp128 (.in0(cmp128_in0), .in1(cmp128_in1), .out0(cmp128_out0), .out1(cmp128_out1));
cmp cmp129 (.in0(cmp129_in0), .in1(cmp129_in1), .out0(cmp129_out0), .out1(cmp129_out1));
cmp cmp130 (.in0(cmp130_in0), .in1(cmp130_in1), .out0(cmp130_out0), .out1(cmp130_out1));
cmp cmp131 (.in0(cmp131_in0), .in1(cmp131_in1), .out0(cmp131_out0), .out1(cmp131_out1));
cmp cmp132 (.in0(cmp132_in0), .in1(cmp132_in1), .out0(cmp132_out0), .out1(cmp132_out1));
cmp cmp133 (.in0(cmp133_in0), .in1(cmp133_in1), .out0(cmp133_out0), .out1(cmp133_out1));
cmp cmp134 (.in0(cmp134_in0), .in1(cmp134_in1), .out0(cmp134_out0), .out1(cmp134_out1));
cmp cmp135 (.in0(cmp135_in0), .in1(cmp135_in1), .out0(cmp135_out0), .out1(cmp135_out1));
cmp cmp136 (.in0(cmp136_in0), .in1(cmp136_in1), .out0(cmp136_out0), .out1(cmp136_out1));
cmp cmp137 (.in0(cmp137_in0), .in1(cmp137_in1), .out0(cmp137_out0), .out1(cmp137_out1));
cmp cmp138 (.in0(cmp138_in0), .in1(cmp138_in1), .out0(cmp138_out0), .out1(cmp138_out1));
cmp cmp139 (.in0(cmp139_in0), .in1(cmp139_in1), .out0(cmp139_out0), .out1(cmp139_out1));
cmp cmp140 (.in0(cmp140_in0), .in1(cmp140_in1), .out0(cmp140_out0), .out1(cmp140_out1));
cmp cmp141 (.in0(cmp141_in0), .in1(cmp141_in1), .out0(cmp141_out0), .out1(cmp141_out1));
cmp cmp142 (.in0(cmp142_in0), .in1(cmp142_in1), .out0(cmp142_out0), .out1(cmp142_out1));
cmp cmp143 (.in0(cmp143_in0), .in1(cmp143_in1), .out0(cmp143_out0), .out1(cmp143_out1));
cmp cmp144 (.in0(cmp144_in0), .in1(cmp144_in1), .out0(cmp144_out0), .out1(cmp144_out1));
cmp cmp145 (.in0(cmp145_in0), .in1(cmp145_in1), .out0(cmp145_out0), .out1(cmp145_out1));
cmp cmp146 (.in0(cmp146_in0), .in1(cmp146_in1), .out0(cmp146_out0), .out1(cmp146_out1));
cmp cmp147 (.in0(cmp147_in0), .in1(cmp147_in1), .out0(cmp147_out0), .out1(cmp147_out1));
cmp cmp148 (.in0(cmp148_in0), .in1(cmp148_in1), .out0(cmp148_out0), .out1(cmp148_out1));
cmp cmp149 (.in0(cmp149_in0), .in1(cmp149_in1), .out0(cmp149_out0), .out1(cmp149_out1));
cmp cmp150 (.in0(cmp150_in0), .in1(cmp150_in1), .out0(cmp150_out0), .out1(cmp150_out1));
cmp cmp151 (.in0(cmp151_in0), .in1(cmp151_in1), .out0(cmp151_out0), .out1(cmp151_out1));
cmp cmp152 (.in0(cmp152_in0), .in1(cmp152_in1), .out0(cmp152_out0), .out1(cmp152_out1));
cmp cmp153 (.in0(cmp153_in0), .in1(cmp153_in1), .out0(cmp153_out0), .out1(cmp153_out1));
cmp cmp154 (.in0(cmp154_in0), .in1(cmp154_in1), .out0(cmp154_out0), .out1(cmp154_out1));
cmp cmp155 (.in0(cmp155_in0), .in1(cmp155_in1), .out0(cmp155_out0), .out1(cmp155_out1));
cmp cmp156 (.in0(cmp156_in0), .in1(cmp156_in1), .out0(cmp156_out0), .out1(cmp156_out1));
cmp cmp157 (.in0(cmp157_in0), .in1(cmp157_in1), .out0(cmp157_out0), .out1(cmp157_out1));
cmp cmp158 (.in0(cmp158_in0), .in1(cmp158_in1), .out0(cmp158_out0), .out1(cmp158_out1));
cmp cmp159 (.in0(cmp159_in0), .in1(cmp159_in1), .out0(cmp159_out0), .out1(cmp159_out1));
cmp cmp160 (.in0(cmp160_in0), .in1(cmp160_in1), .out0(cmp160_out0), .out1(cmp160_out1));
cmp cmp161 (.in0(cmp161_in0), .in1(cmp161_in1), .out0(cmp161_out0), .out1(cmp161_out1));
cmp cmp162 (.in0(cmp162_in0), .in1(cmp162_in1), .out0(cmp162_out0), .out1(cmp162_out1));
cmp cmp163 (.in0(cmp163_in0), .in1(cmp163_in1), .out0(cmp163_out0), .out1(cmp163_out1));
cmp cmp164 (.in0(cmp164_in0), .in1(cmp164_in1), .out0(cmp164_out0), .out1(cmp164_out1));
cmp cmp165 (.in0(cmp165_in0), .in1(cmp165_in1), .out0(cmp165_out0), .out1(cmp165_out1));
cmp cmp166 (.in0(cmp166_in0), .in1(cmp166_in1), .out0(cmp166_out0), .out1(cmp166_out1));
cmp cmp167 (.in0(cmp167_in0), .in1(cmp167_in1), .out0(cmp167_out0), .out1(cmp167_out1));
cmp cmp168 (.in0(cmp168_in0), .in1(cmp168_in1), .out0(cmp168_out0), .out1(cmp168_out1));
cmp cmp169 (.in0(cmp169_in0), .in1(cmp169_in1), .out0(cmp169_out0), .out1(cmp169_out1));
cmp cmp170 (.in0(cmp170_in0), .in1(cmp170_in1), .out0(cmp170_out0), .out1(cmp170_out1));
cmp cmp171 (.in0(cmp171_in0), .in1(cmp171_in1), .out0(cmp171_out0), .out1(cmp171_out1));
cmp cmp172 (.in0(cmp172_in0), .in1(cmp172_in1), .out0(cmp172_out0), .out1(cmp172_out1));
cmp cmp173 (.in0(cmp173_in0), .in1(cmp173_in1), .out0(cmp173_out0), .out1(cmp173_out1));
cmp cmp174 (.in0(cmp174_in0), .in1(cmp174_in1), .out0(cmp174_out0), .out1(cmp174_out1));
cmp cmp175 (.in0(cmp175_in0), .in1(cmp175_in1), .out0(cmp175_out0), .out1(cmp175_out1));
cmp cmp176 (.in0(cmp176_in0), .in1(cmp176_in1), .out0(cmp176_out0), .out1(cmp176_out1));
cmp cmp177 (.in0(cmp177_in0), .in1(cmp177_in1), .out0(cmp177_out0), .out1(cmp177_out1));
cmp cmp178 (.in0(cmp178_in0), .in1(cmp178_in1), .out0(cmp178_out0), .out1(cmp178_out1));
cmp cmp179 (.in0(cmp179_in0), .in1(cmp179_in1), .out0(cmp179_out0), .out1(cmp179_out1));
cmp cmp180 (.in0(cmp180_in0), .in1(cmp180_in1), .out0(cmp180_out0), .out1(cmp180_out1));
cmp cmp181 (.in0(cmp181_in0), .in1(cmp181_in1), .out0(cmp181_out0), .out1(cmp181_out1));
cmp cmp182 (.in0(cmp182_in0), .in1(cmp182_in1), .out0(cmp182_out0), .out1(cmp182_out1));
cmp cmp183 (.in0(cmp183_in0), .in1(cmp183_in1), .out0(cmp183_out0), .out1(cmp183_out1));
cmp cmp184 (.in0(cmp184_in0), .in1(cmp184_in1), .out0(cmp184_out0), .out1(cmp184_out1));
cmp cmp185 (.in0(cmp185_in0), .in1(cmp185_in1), .out0(cmp185_out0), .out1(cmp185_out1));
cmp cmp186 (.in0(cmp186_in0), .in1(cmp186_in1), .out0(cmp186_out0), .out1(cmp186_out1));
cmp cmp187 (.in0(cmp187_in0), .in1(cmp187_in1), .out0(cmp187_out0), .out1(cmp187_out1));
cmp cmp188 (.in0(cmp188_in0), .in1(cmp188_in1), .out0(cmp188_out0), .out1(cmp188_out1));
cmp cmp189 (.in0(cmp189_in0), .in1(cmp189_in1), .out0(cmp189_out0), .out1(cmp189_out1));
cmp cmp190 (.in0(cmp190_in0), .in1(cmp190_in1), .out0(cmp190_out0), .out1(cmp190_out1));
cmp cmp191 (.in0(cmp191_in0), .in1(cmp191_in1), .out0(cmp191_out0), .out1(cmp191_out1));
cmp cmp192 (.in0(cmp192_in0), .in1(cmp192_in1), .out0(cmp192_out0), .out1(cmp192_out1));
cmp cmp193 (.in0(cmp193_in0), .in1(cmp193_in1), .out0(cmp193_out0), .out1(cmp193_out1));
cmp cmp194 (.in0(cmp194_in0), .in1(cmp194_in1), .out0(cmp194_out0), .out1(cmp194_out1));
cmp cmp195 (.in0(cmp195_in0), .in1(cmp195_in1), .out0(cmp195_out0), .out1(cmp195_out1));
cmp cmp196 (.in0(cmp196_in0), .in1(cmp196_in1), .out0(cmp196_out0), .out1(cmp196_out1));
cmp cmp197 (.in0(cmp197_in0), .in1(cmp197_in1), .out0(cmp197_out0), .out1(cmp197_out1));
cmp cmp198 (.in0(cmp198_in0), .in1(cmp198_in1), .out0(cmp198_out0), .out1(cmp198_out1));
cmp cmp199 (.in0(cmp199_in0), .in1(cmp199_in1), .out0(cmp199_out0), .out1(cmp199_out1));
cmp cmp200 (.in0(cmp200_in0), .in1(cmp200_in1), .out0(cmp200_out0), .out1(cmp200_out1));
cmp cmp201 (.in0(cmp201_in0), .in1(cmp201_in1), .out0(cmp201_out0), .out1(cmp201_out1));
cmp cmp202 (.in0(cmp202_in0), .in1(cmp202_in1), .out0(cmp202_out0), .out1(cmp202_out1));
cmp cmp203 (.in0(cmp203_in0), .in1(cmp203_in1), .out0(cmp203_out0), .out1(cmp203_out1));
cmp cmp204 (.in0(cmp204_in0), .in1(cmp204_in1), .out0(cmp204_out0), .out1(cmp204_out1));
cmp cmp205 (.in0(cmp205_in0), .in1(cmp205_in1), .out0(cmp205_out0), .out1(cmp205_out1));
cmp cmp206 (.in0(cmp206_in0), .in1(cmp206_in1), .out0(cmp206_out0), .out1(cmp206_out1));
cmp cmp207 (.in0(cmp207_in0), .in1(cmp207_in1), .out0(cmp207_out0), .out1(cmp207_out1));
cmp cmp208 (.in0(cmp208_in0), .in1(cmp208_in1), .out0(cmp208_out0), .out1(cmp208_out1));
cmp cmp209 (.in0(cmp209_in0), .in1(cmp209_in1), .out0(cmp209_out0), .out1(cmp209_out1));
cmp cmp210 (.in0(cmp210_in0), .in1(cmp210_in1), .out0(cmp210_out0), .out1(cmp210_out1));
cmp cmp211 (.in0(cmp211_in0), .in1(cmp211_in1), .out0(cmp211_out0), .out1(cmp211_out1));
cmp cmp212 (.in0(cmp212_in0), .in1(cmp212_in1), .out0(cmp212_out0), .out1(cmp212_out1));
cmp cmp213 (.in0(cmp213_in0), .in1(cmp213_in1), .out0(cmp213_out0), .out1(cmp213_out1));
cmp cmp214 (.in0(cmp214_in0), .in1(cmp214_in1), .out0(cmp214_out0), .out1(cmp214_out1));
cmp cmp215 (.in0(cmp215_in0), .in1(cmp215_in1), .out0(cmp215_out0), .out1(cmp215_out1));
cmp cmp216 (.in0(cmp216_in0), .in1(cmp216_in1), .out0(cmp216_out0), .out1(cmp216_out1));
cmp cmp217 (.in0(cmp217_in0), .in1(cmp217_in1), .out0(cmp217_out0), .out1(cmp217_out1));
cmp cmp218 (.in0(cmp218_in0), .in1(cmp218_in1), .out0(cmp218_out0), .out1(cmp218_out1));
cmp cmp219 (.in0(cmp219_in0), .in1(cmp219_in1), .out0(cmp219_out0), .out1(cmp219_out1));
cmp cmp220 (.in0(cmp220_in0), .in1(cmp220_in1), .out0(cmp220_out0), .out1(cmp220_out1));
cmp cmp221 (.in0(cmp221_in0), .in1(cmp221_in1), .out0(cmp221_out0), .out1(cmp221_out1));
cmp cmp222 (.in0(cmp222_in0), .in1(cmp222_in1), .out0(cmp222_out0), .out1(cmp222_out1));
cmp cmp223 (.in0(cmp223_in0), .in1(cmp223_in1), .out0(cmp223_out0), .out1(cmp223_out1));
cmp cmp224 (.in0(cmp224_in0), .in1(cmp224_in1), .out0(cmp224_out0), .out1(cmp224_out1));
cmp cmp225 (.in0(cmp225_in0), .in1(cmp225_in1), .out0(cmp225_out0), .out1(cmp225_out1));
cmp cmp226 (.in0(cmp226_in0), .in1(cmp226_in1), .out0(cmp226_out0), .out1(cmp226_out1));
cmp cmp227 (.in0(cmp227_in0), .in1(cmp227_in1), .out0(cmp227_out0), .out1(cmp227_out1));
cmp cmp228 (.in0(cmp228_in0), .in1(cmp228_in1), .out0(cmp228_out0), .out1(cmp228_out1));
cmp cmp229 (.in0(cmp229_in0), .in1(cmp229_in1), .out0(cmp229_out0), .out1(cmp229_out1));
cmp cmp230 (.in0(cmp230_in0), .in1(cmp230_in1), .out0(cmp230_out0), .out1(cmp230_out1));
cmp cmp231 (.in0(cmp231_in0), .in1(cmp231_in1), .out0(cmp231_out0), .out1(cmp231_out1));
cmp cmp232 (.in0(cmp232_in0), .in1(cmp232_in1), .out0(cmp232_out0), .out1(cmp232_out1));
cmp cmp233 (.in0(cmp233_in0), .in1(cmp233_in1), .out0(cmp233_out0), .out1(cmp233_out1));
cmp cmp234 (.in0(cmp234_in0), .in1(cmp234_in1), .out0(cmp234_out0), .out1(cmp234_out1));
cmp cmp235 (.in0(cmp235_in0), .in1(cmp235_in1), .out0(cmp235_out0), .out1(cmp235_out1));
cmp cmp236 (.in0(cmp236_in0), .in1(cmp236_in1), .out0(cmp236_out0), .out1(cmp236_out1));
cmp cmp237 (.in0(cmp237_in0), .in1(cmp237_in1), .out0(cmp237_out0), .out1(cmp237_out1));
cmp cmp238 (.in0(cmp238_in0), .in1(cmp238_in1), .out0(cmp238_out0), .out1(cmp238_out1));
cmp cmp239 (.in0(cmp239_in0), .in1(cmp239_in1), .out0(cmp239_out0), .out1(cmp239_out1));
cmp cmp240 (.in0(cmp240_in0), .in1(cmp240_in1), .out0(cmp240_out0), .out1(cmp240_out1));
cmp cmp241 (.in0(cmp241_in0), .in1(cmp241_in1), .out0(cmp241_out0), .out1(cmp241_out1));
cmp cmp242 (.in0(cmp242_in0), .in1(cmp242_in1), .out0(cmp242_out0), .out1(cmp242_out1));
cmp cmp243 (.in0(cmp243_in0), .in1(cmp243_in1), .out0(cmp243_out0), .out1(cmp243_out1));
cmp cmp244 (.in0(cmp244_in0), .in1(cmp244_in1), .out0(cmp244_out0), .out1(cmp244_out1));
cmp cmp245 (.in0(cmp245_in0), .in1(cmp245_in1), .out0(cmp245_out0), .out1(cmp245_out1));
cmp cmp246 (.in0(cmp246_in0), .in1(cmp246_in1), .out0(cmp246_out0), .out1(cmp246_out1));
cmp cmp247 (.in0(cmp247_in0), .in1(cmp247_in1), .out0(cmp247_out0), .out1(cmp247_out1));
cmp cmp248 (.in0(cmp248_in0), .in1(cmp248_in1), .out0(cmp248_out0), .out1(cmp248_out1));
cmp cmp249 (.in0(cmp249_in0), .in1(cmp249_in1), .out0(cmp249_out0), .out1(cmp249_out1));
cmp cmp250 (.in0(cmp250_in0), .in1(cmp250_in1), .out0(cmp250_out0), .out1(cmp250_out1));
cmp cmp251 (.in0(cmp251_in0), .in1(cmp251_in1), .out0(cmp251_out0), .out1(cmp251_out1));
cmp cmp252 (.in0(cmp252_in0), .in1(cmp252_in1), .out0(cmp252_out0), .out1(cmp252_out1));
cmp cmp253 (.in0(cmp253_in0), .in1(cmp253_in1), .out0(cmp253_out0), .out1(cmp253_out1));
cmp cmp254 (.in0(cmp254_in0), .in1(cmp254_in1), .out0(cmp254_out0), .out1(cmp254_out1));
cmp cmp255 (.in0(cmp255_in0), .in1(cmp255_in1), .out0(cmp255_out0), .out1(cmp255_out1));
cmp cmp256 (.in0(cmp256_in0), .in1(cmp256_in1), .out0(cmp256_out0), .out1(cmp256_out1));
cmp cmp257 (.in0(cmp257_in0), .in1(cmp257_in1), .out0(cmp257_out0), .out1(cmp257_out1));
cmp cmp258 (.in0(cmp258_in0), .in1(cmp258_in1), .out0(cmp258_out0), .out1(cmp258_out1));
cmp cmp259 (.in0(cmp259_in0), .in1(cmp259_in1), .out0(cmp259_out0), .out1(cmp259_out1));
cmp cmp260 (.in0(cmp260_in0), .in1(cmp260_in1), .out0(cmp260_out0), .out1(cmp260_out1));
cmp cmp261 (.in0(cmp261_in0), .in1(cmp261_in1), .out0(cmp261_out0), .out1(cmp261_out1));
cmp cmp262 (.in0(cmp262_in0), .in1(cmp262_in1), .out0(cmp262_out0), .out1(cmp262_out1));
cmp cmp263 (.in0(cmp263_in0), .in1(cmp263_in1), .out0(cmp263_out0), .out1(cmp263_out1));
cmp cmp264 (.in0(cmp264_in0), .in1(cmp264_in1), .out0(cmp264_out0), .out1(cmp264_out1));
cmp cmp265 (.in0(cmp265_in0), .in1(cmp265_in1), .out0(cmp265_out0), .out1(cmp265_out1));
cmp cmp266 (.in0(cmp266_in0), .in1(cmp266_in1), .out0(cmp266_out0), .out1(cmp266_out1));
cmp cmp267 (.in0(cmp267_in0), .in1(cmp267_in1), .out0(cmp267_out0), .out1(cmp267_out1));
cmp cmp268 (.in0(cmp268_in0), .in1(cmp268_in1), .out0(cmp268_out0), .out1(cmp268_out1));
cmp cmp269 (.in0(cmp269_in0), .in1(cmp269_in1), .out0(cmp269_out0), .out1(cmp269_out1));
cmp cmp270 (.in0(cmp270_in0), .in1(cmp270_in1), .out0(cmp270_out0), .out1(cmp270_out1));
cmp cmp271 (.in0(cmp271_in0), .in1(cmp271_in1), .out0(cmp271_out0), .out1(cmp271_out1));
cmp cmp272 (.in0(cmp272_in0), .in1(cmp272_in1), .out0(cmp272_out0), .out1(cmp272_out1));
cmp cmp273 (.in0(cmp273_in0), .in1(cmp273_in1), .out0(cmp273_out0), .out1(cmp273_out1));
cmp cmp274 (.in0(cmp274_in0), .in1(cmp274_in1), .out0(cmp274_out0), .out1(cmp274_out1));
cmp cmp275 (.in0(cmp275_in0), .in1(cmp275_in1), .out0(cmp275_out0), .out1(cmp275_out1));
cmp cmp276 (.in0(cmp276_in0), .in1(cmp276_in1), .out0(cmp276_out0), .out1(cmp276_out1));
cmp cmp277 (.in0(cmp277_in0), .in1(cmp277_in1), .out0(cmp277_out0), .out1(cmp277_out1));
cmp cmp278 (.in0(cmp278_in0), .in1(cmp278_in1), .out0(cmp278_out0), .out1(cmp278_out1));
cmp cmp279 (.in0(cmp279_in0), .in1(cmp279_in1), .out0(cmp279_out0), .out1(cmp279_out1));
cmp cmp280 (.in0(cmp280_in0), .in1(cmp280_in1), .out0(cmp280_out0), .out1(cmp280_out1));
cmp cmp281 (.in0(cmp281_in0), .in1(cmp281_in1), .out0(cmp281_out0), .out1(cmp281_out1));
cmp cmp282 (.in0(cmp282_in0), .in1(cmp282_in1), .out0(cmp282_out0), .out1(cmp282_out1));
cmp cmp283 (.in0(cmp283_in0), .in1(cmp283_in1), .out0(cmp283_out0), .out1(cmp283_out1));
cmp cmp284 (.in0(cmp284_in0), .in1(cmp284_in1), .out0(cmp284_out0), .out1(cmp284_out1));
cmp cmp285 (.in0(cmp285_in0), .in1(cmp285_in1), .out0(cmp285_out0), .out1(cmp285_out1));
cmp cmp286 (.in0(cmp286_in0), .in1(cmp286_in1), .out0(cmp286_out0), .out1(cmp286_out1));
cmp cmp287 (.in0(cmp287_in0), .in1(cmp287_in1), .out0(cmp287_out0), .out1(cmp287_out1));
cmp cmp288 (.in0(cmp288_in0), .in1(cmp288_in1), .out0(cmp288_out0), .out1(cmp288_out1));
cmp cmp289 (.in0(cmp289_in0), .in1(cmp289_in1), .out0(cmp289_out0), .out1(cmp289_out1));
cmp cmp290 (.in0(cmp290_in0), .in1(cmp290_in1), .out0(cmp290_out0), .out1(cmp290_out1));
cmp cmp291 (.in0(cmp291_in0), .in1(cmp291_in1), .out0(cmp291_out0), .out1(cmp291_out1));
cmp cmp292 (.in0(cmp292_in0), .in1(cmp292_in1), .out0(cmp292_out0), .out1(cmp292_out1));
cmp cmp293 (.in0(cmp293_in0), .in1(cmp293_in1), .out0(cmp293_out0), .out1(cmp293_out1));
cmp cmp294 (.in0(cmp294_in0), .in1(cmp294_in1), .out0(cmp294_out0), .out1(cmp294_out1));
cmp cmp295 (.in0(cmp295_in0), .in1(cmp295_in1), .out0(cmp295_out0), .out1(cmp295_out1));
cmp cmp296 (.in0(cmp296_in0), .in1(cmp296_in1), .out0(cmp296_out0), .out1(cmp296_out1));
cmp cmp297 (.in0(cmp297_in0), .in1(cmp297_in1), .out0(cmp297_out0), .out1(cmp297_out1));
cmp cmp298 (.in0(cmp298_in0), .in1(cmp298_in1), .out0(cmp298_out0), .out1(cmp298_out1));
cmp cmp299 (.in0(cmp299_in0), .in1(cmp299_in1), .out0(cmp299_out0), .out1(cmp299_out1));
cmp cmp300 (.in0(cmp300_in0), .in1(cmp300_in1), .out0(cmp300_out0), .out1(cmp300_out1));
cmp cmp301 (.in0(cmp301_in0), .in1(cmp301_in1), .out0(cmp301_out0), .out1(cmp301_out1));
cmp cmp302 (.in0(cmp302_in0), .in1(cmp302_in1), .out0(cmp302_out0), .out1(cmp302_out1));
cmp cmp303 (.in0(cmp303_in0), .in1(cmp303_in1), .out0(cmp303_out0), .out1(cmp303_out1));
cmp cmp304 (.in0(cmp304_in0), .in1(cmp304_in1), .out0(cmp304_out0), .out1(cmp304_out1));
cmp cmp305 (.in0(cmp305_in0), .in1(cmp305_in1), .out0(cmp305_out0), .out1(cmp305_out1));
cmp cmp306 (.in0(cmp306_in0), .in1(cmp306_in1), .out0(cmp306_out0), .out1(cmp306_out1));
cmp cmp307 (.in0(cmp307_in0), .in1(cmp307_in1), .out0(cmp307_out0), .out1(cmp307_out1));
cmp cmp308 (.in0(cmp308_in0), .in1(cmp308_in1), .out0(cmp308_out0), .out1(cmp308_out1));
cmp cmp309 (.in0(cmp309_in0), .in1(cmp309_in1), .out0(cmp309_out0), .out1(cmp309_out1));
cmp cmp310 (.in0(cmp310_in0), .in1(cmp310_in1), .out0(cmp310_out0), .out1(cmp310_out1));
cmp cmp311 (.in0(cmp311_in0), .in1(cmp311_in1), .out0(cmp311_out0), .out1(cmp311_out1));
cmp cmp312 (.in0(cmp312_in0), .in1(cmp312_in1), .out0(cmp312_out0), .out1(cmp312_out1));
cmp cmp313 (.in0(cmp313_in0), .in1(cmp313_in1), .out0(cmp313_out0), .out1(cmp313_out1));
cmp cmp314 (.in0(cmp314_in0), .in1(cmp314_in1), .out0(cmp314_out0), .out1(cmp314_out1));
cmp cmp315 (.in0(cmp315_in0), .in1(cmp315_in1), .out0(cmp315_out0), .out1(cmp315_out1));
cmp cmp316 (.in0(cmp316_in0), .in1(cmp316_in1), .out0(cmp316_out0), .out1(cmp316_out1));
cmp cmp317 (.in0(cmp317_in0), .in1(cmp317_in1), .out0(cmp317_out0), .out1(cmp317_out1));
cmp cmp318 (.in0(cmp318_in0), .in1(cmp318_in1), .out0(cmp318_out0), .out1(cmp318_out1));
cmp cmp319 (.in0(cmp319_in0), .in1(cmp319_in1), .out0(cmp319_out0), .out1(cmp319_out1));
cmp cmp320 (.in0(cmp320_in0), .in1(cmp320_in1), .out0(cmp320_out0), .out1(cmp320_out1));
cmp cmp321 (.in0(cmp321_in0), .in1(cmp321_in1), .out0(cmp321_out0), .out1(cmp321_out1));
cmp cmp322 (.in0(cmp322_in0), .in1(cmp322_in1), .out0(cmp322_out0), .out1(cmp322_out1));
cmp cmp323 (.in0(cmp323_in0), .in1(cmp323_in1), .out0(cmp323_out0), .out1(cmp323_out1));
cmp cmp324 (.in0(cmp324_in0), .in1(cmp324_in1), .out0(cmp324_out0), .out1(cmp324_out1));
cmp cmp325 (.in0(cmp325_in0), .in1(cmp325_in1), .out0(cmp325_out0), .out1(cmp325_out1));
cmp cmp326 (.in0(cmp326_in0), .in1(cmp326_in1), .out0(cmp326_out0), .out1(cmp326_out1));
cmp cmp327 (.in0(cmp327_in0), .in1(cmp327_in1), .out0(cmp327_out0), .out1(cmp327_out1));
cmp cmp328 (.in0(cmp328_in0), .in1(cmp328_in1), .out0(cmp328_out0), .out1(cmp328_out1));
cmp cmp329 (.in0(cmp329_in0), .in1(cmp329_in1), .out0(cmp329_out0), .out1(cmp329_out1));
cmp cmp330 (.in0(cmp330_in0), .in1(cmp330_in1), .out0(cmp330_out0), .out1(cmp330_out1));
cmp cmp331 (.in0(cmp331_in0), .in1(cmp331_in1), .out0(cmp331_out0), .out1(cmp331_out1));
cmp cmp332 (.in0(cmp332_in0), .in1(cmp332_in1), .out0(cmp332_out0), .out1(cmp332_out1));
cmp cmp333 (.in0(cmp333_in0), .in1(cmp333_in1), .out0(cmp333_out0), .out1(cmp333_out1));
cmp cmp334 (.in0(cmp334_in0), .in1(cmp334_in1), .out0(cmp334_out0), .out1(cmp334_out1));
cmp cmp335 (.in0(cmp335_in0), .in1(cmp335_in1), .out0(cmp335_out0), .out1(cmp335_out1));
cmp cmp336 (.in0(cmp336_in0), .in1(cmp336_in1), .out0(cmp336_out0), .out1(cmp336_out1));
cmp cmp337 (.in0(cmp337_in0), .in1(cmp337_in1), .out0(cmp337_out0), .out1(cmp337_out1));
cmp cmp338 (.in0(cmp338_in0), .in1(cmp338_in1), .out0(cmp338_out0), .out1(cmp338_out1));
cmp cmp339 (.in0(cmp339_in0), .in1(cmp339_in1), .out0(cmp339_out0), .out1(cmp339_out1));
cmp cmp340 (.in0(cmp340_in0), .in1(cmp340_in1), .out0(cmp340_out0), .out1(cmp340_out1));
cmp cmp341 (.in0(cmp341_in0), .in1(cmp341_in1), .out0(cmp341_out0), .out1(cmp341_out1));
cmp cmp342 (.in0(cmp342_in0), .in1(cmp342_in1), .out0(cmp342_out0), .out1(cmp342_out1));
cmp cmp343 (.in0(cmp343_in0), .in1(cmp343_in1), .out0(cmp343_out0), .out1(cmp343_out1));
cmp cmp344 (.in0(cmp344_in0), .in1(cmp344_in1), .out0(cmp344_out0), .out1(cmp344_out1));
cmp cmp345 (.in0(cmp345_in0), .in1(cmp345_in1), .out0(cmp345_out0), .out1(cmp345_out1));
cmp cmp346 (.in0(cmp346_in0), .in1(cmp346_in1), .out0(cmp346_out0), .out1(cmp346_out1));
cmp cmp347 (.in0(cmp347_in0), .in1(cmp347_in1), .out0(cmp347_out0), .out1(cmp347_out1));
cmp cmp348 (.in0(cmp348_in0), .in1(cmp348_in1), .out0(cmp348_out0), .out1(cmp348_out1));
cmp cmp349 (.in0(cmp349_in0), .in1(cmp349_in1), .out0(cmp349_out0), .out1(cmp349_out1));
cmp cmp350 (.in0(cmp350_in0), .in1(cmp350_in1), .out0(cmp350_out0), .out1(cmp350_out1));
cmp cmp351 (.in0(cmp351_in0), .in1(cmp351_in1), .out0(cmp351_out0), .out1(cmp351_out1));
cmp cmp352 (.in0(cmp352_in0), .in1(cmp352_in1), .out0(cmp352_out0), .out1(cmp352_out1));
cmp cmp353 (.in0(cmp353_in0), .in1(cmp353_in1), .out0(cmp353_out0), .out1(cmp353_out1));
cmp cmp354 (.in0(cmp354_in0), .in1(cmp354_in1), .out0(cmp354_out0), .out1(cmp354_out1));
cmp cmp355 (.in0(cmp355_in0), .in1(cmp355_in1), .out0(cmp355_out0), .out1(cmp355_out1));
cmp cmp356 (.in0(cmp356_in0), .in1(cmp356_in1), .out0(cmp356_out0), .out1(cmp356_out1));
cmp cmp357 (.in0(cmp357_in0), .in1(cmp357_in1), .out0(cmp357_out0), .out1(cmp357_out1));
cmp cmp358 (.in0(cmp358_in0), .in1(cmp358_in1), .out0(cmp358_out0), .out1(cmp358_out1));
cmp cmp359 (.in0(cmp359_in0), .in1(cmp359_in1), .out0(cmp359_out0), .out1(cmp359_out1));
cmp cmp360 (.in0(cmp360_in0), .in1(cmp360_in1), .out0(cmp360_out0), .out1(cmp360_out1));
cmp cmp361 (.in0(cmp361_in0), .in1(cmp361_in1), .out0(cmp361_out0), .out1(cmp361_out1));
cmp cmp362 (.in0(cmp362_in0), .in1(cmp362_in1), .out0(cmp362_out0), .out1(cmp362_out1));
cmp cmp363 (.in0(cmp363_in0), .in1(cmp363_in1), .out0(cmp363_out0), .out1(cmp363_out1));
cmp cmp364 (.in0(cmp364_in0), .in1(cmp364_in1), .out0(cmp364_out0), .out1(cmp364_out1));
cmp cmp365 (.in0(cmp365_in0), .in1(cmp365_in1), .out0(cmp365_out0), .out1(cmp365_out1));
cmp cmp366 (.in0(cmp366_in0), .in1(cmp366_in1), .out0(cmp366_out0), .out1(cmp366_out1));
cmp cmp367 (.in0(cmp367_in0), .in1(cmp367_in1), .out0(cmp367_out0), .out1(cmp367_out1));
cmp cmp368 (.in0(cmp368_in0), .in1(cmp368_in1), .out0(cmp368_out0), .out1(cmp368_out1));
cmp cmp369 (.in0(cmp369_in0), .in1(cmp369_in1), .out0(cmp369_out0), .out1(cmp369_out1));
cmp cmp370 (.in0(cmp370_in0), .in1(cmp370_in1), .out0(cmp370_out0), .out1(cmp370_out1));
cmp cmp371 (.in0(cmp371_in0), .in1(cmp371_in1), .out0(cmp371_out0), .out1(cmp371_out1));
cmp cmp372 (.in0(cmp372_in0), .in1(cmp372_in1), .out0(cmp372_out0), .out1(cmp372_out1));
cmp cmp373 (.in0(cmp373_in0), .in1(cmp373_in1), .out0(cmp373_out0), .out1(cmp373_out1));
cmp cmp374 (.in0(cmp374_in0), .in1(cmp374_in1), .out0(cmp374_out0), .out1(cmp374_out1));
cmp cmp375 (.in0(cmp375_in0), .in1(cmp375_in1), .out0(cmp375_out0), .out1(cmp375_out1));
cmp cmp376 (.in0(cmp376_in0), .in1(cmp376_in1), .out0(cmp376_out0), .out1(cmp376_out1));
cmp cmp377 (.in0(cmp377_in0), .in1(cmp377_in1), .out0(cmp377_out0), .out1(cmp377_out1));
cmp cmp378 (.in0(cmp378_in0), .in1(cmp378_in1), .out0(cmp378_out0), .out1(cmp378_out1));
cmp cmp379 (.in0(cmp379_in0), .in1(cmp379_in1), .out0(cmp379_out0), .out1(cmp379_out1));
cmp cmp380 (.in0(cmp380_in0), .in1(cmp380_in1), .out0(cmp380_out0), .out1(cmp380_out1));
cmp cmp381 (.in0(cmp381_in0), .in1(cmp381_in1), .out0(cmp381_out0), .out1(cmp381_out1));
cmp cmp382 (.in0(cmp382_in0), .in1(cmp382_in1), .out0(cmp382_out0), .out1(cmp382_out1));
cmp cmp383 (.in0(cmp383_in0), .in1(cmp383_in1), .out0(cmp383_out0), .out1(cmp383_out1));
cmp cmp384 (.in0(cmp384_in0), .in1(cmp384_in1), .out0(cmp384_out0), .out1(cmp384_out1));
cmp cmp385 (.in0(cmp385_in0), .in1(cmp385_in1), .out0(cmp385_out0), .out1(cmp385_out1));
cmp cmp386 (.in0(cmp386_in0), .in1(cmp386_in1), .out0(cmp386_out0), .out1(cmp386_out1));
cmp cmp387 (.in0(cmp387_in0), .in1(cmp387_in1), .out0(cmp387_out0), .out1(cmp387_out1));
cmp cmp388 (.in0(cmp388_in0), .in1(cmp388_in1), .out0(cmp388_out0), .out1(cmp388_out1));
cmp cmp389 (.in0(cmp389_in0), .in1(cmp389_in1), .out0(cmp389_out0), .out1(cmp389_out1));
cmp cmp390 (.in0(cmp390_in0), .in1(cmp390_in1), .out0(cmp390_out0), .out1(cmp390_out1));
cmp cmp391 (.in0(cmp391_in0), .in1(cmp391_in1), .out0(cmp391_out0), .out1(cmp391_out1));
cmp cmp392 (.in0(cmp392_in0), .in1(cmp392_in1), .out0(cmp392_out0), .out1(cmp392_out1));
cmp cmp393 (.in0(cmp393_in0), .in1(cmp393_in1), .out0(cmp393_out0), .out1(cmp393_out1));
cmp cmp394 (.in0(cmp394_in0), .in1(cmp394_in1), .out0(cmp394_out0), .out1(cmp394_out1));
cmp cmp395 (.in0(cmp395_in0), .in1(cmp395_in1), .out0(cmp395_out0), .out1(cmp395_out1));
cmp cmp396 (.in0(cmp396_in0), .in1(cmp396_in1), .out0(cmp396_out0), .out1(cmp396_out1));
cmp cmp397 (.in0(cmp397_in0), .in1(cmp397_in1), .out0(cmp397_out0), .out1(cmp397_out1));
cmp cmp398 (.in0(cmp398_in0), .in1(cmp398_in1), .out0(cmp398_out0), .out1(cmp398_out1));
cmp cmp399 (.in0(cmp399_in0), .in1(cmp399_in1), .out0(cmp399_out0), .out1(cmp399_out1));
cmp cmp400 (.in0(cmp400_in0), .in1(cmp400_in1), .out0(cmp400_out0), .out1(cmp400_out1));
cmp cmp401 (.in0(cmp401_in0), .in1(cmp401_in1), .out0(cmp401_out0), .out1(cmp401_out1));
cmp cmp402 (.in0(cmp402_in0), .in1(cmp402_in1), .out0(cmp402_out0), .out1(cmp402_out1));
cmp cmp403 (.in0(cmp403_in0), .in1(cmp403_in1), .out0(cmp403_out0), .out1(cmp403_out1));
cmp cmp404 (.in0(cmp404_in0), .in1(cmp404_in1), .out0(cmp404_out0), .out1(cmp404_out1));
cmp cmp405 (.in0(cmp405_in0), .in1(cmp405_in1), .out0(cmp405_out0), .out1(cmp405_out1));
cmp cmp406 (.in0(cmp406_in0), .in1(cmp406_in1), .out0(cmp406_out0), .out1(cmp406_out1));
cmp cmp407 (.in0(cmp407_in0), .in1(cmp407_in1), .out0(cmp407_out0), .out1(cmp407_out1));
cmp cmp408 (.in0(cmp408_in0), .in1(cmp408_in1), .out0(cmp408_out0), .out1(cmp408_out1));
cmp cmp409 (.in0(cmp409_in0), .in1(cmp409_in1), .out0(cmp409_out0), .out1(cmp409_out1));
cmp cmp410 (.in0(cmp410_in0), .in1(cmp410_in1), .out0(cmp410_out0), .out1(cmp410_out1));
cmp cmp411 (.in0(cmp411_in0), .in1(cmp411_in1), .out0(cmp411_out0), .out1(cmp411_out1));
cmp cmp412 (.in0(cmp412_in0), .in1(cmp412_in1), .out0(cmp412_out0), .out1(cmp412_out1));
cmp cmp413 (.in0(cmp413_in0), .in1(cmp413_in1), .out0(cmp413_out0), .out1(cmp413_out1));
cmp cmp414 (.in0(cmp414_in0), .in1(cmp414_in1), .out0(cmp414_out0), .out1(cmp414_out1));
cmp cmp415 (.in0(cmp415_in0), .in1(cmp415_in1), .out0(cmp415_out0), .out1(cmp415_out1));
cmp cmp416 (.in0(cmp416_in0), .in1(cmp416_in1), .out0(cmp416_out0), .out1(cmp416_out1));
cmp cmp417 (.in0(cmp417_in0), .in1(cmp417_in1), .out0(cmp417_out0), .out1(cmp417_out1));
cmp cmp418 (.in0(cmp418_in0), .in1(cmp418_in1), .out0(cmp418_out0), .out1(cmp418_out1));
cmp cmp419 (.in0(cmp419_in0), .in1(cmp419_in1), .out0(cmp419_out0), .out1(cmp419_out1));
cmp cmp420 (.in0(cmp420_in0), .in1(cmp420_in1), .out0(cmp420_out0), .out1(cmp420_out1));
cmp cmp421 (.in0(cmp421_in0), .in1(cmp421_in1), .out0(cmp421_out0), .out1(cmp421_out1));
cmp cmp422 (.in0(cmp422_in0), .in1(cmp422_in1), .out0(cmp422_out0), .out1(cmp422_out1));
cmp cmp423 (.in0(cmp423_in0), .in1(cmp423_in1), .out0(cmp423_out0), .out1(cmp423_out1));
cmp cmp424 (.in0(cmp424_in0), .in1(cmp424_in1), .out0(cmp424_out0), .out1(cmp424_out1));
cmp cmp425 (.in0(cmp425_in0), .in1(cmp425_in1), .out0(cmp425_out0), .out1(cmp425_out1));
cmp cmp426 (.in0(cmp426_in0), .in1(cmp426_in1), .out0(cmp426_out0), .out1(cmp426_out1));
cmp cmp427 (.in0(cmp427_in0), .in1(cmp427_in1), .out0(cmp427_out0), .out1(cmp427_out1));
cmp cmp428 (.in0(cmp428_in0), .in1(cmp428_in1), .out0(cmp428_out0), .out1(cmp428_out1));
cmp cmp429 (.in0(cmp429_in0), .in1(cmp429_in1), .out0(cmp429_out0), .out1(cmp429_out1));
cmp cmp430 (.in0(cmp430_in0), .in1(cmp430_in1), .out0(cmp430_out0), .out1(cmp430_out1));
cmp cmp431 (.in0(cmp431_in0), .in1(cmp431_in1), .out0(cmp431_out0), .out1(cmp431_out1));
cmp cmp432 (.in0(cmp432_in0), .in1(cmp432_in1), .out0(cmp432_out0), .out1(cmp432_out1));
cmp cmp433 (.in0(cmp433_in0), .in1(cmp433_in1), .out0(cmp433_out0), .out1(cmp433_out1));
cmp cmp434 (.in0(cmp434_in0), .in1(cmp434_in1), .out0(cmp434_out0), .out1(cmp434_out1));
cmp cmp435 (.in0(cmp435_in0), .in1(cmp435_in1), .out0(cmp435_out0), .out1(cmp435_out1));
cmp cmp436 (.in0(cmp436_in0), .in1(cmp436_in1), .out0(cmp436_out0), .out1(cmp436_out1));
cmp cmp437 (.in0(cmp437_in0), .in1(cmp437_in1), .out0(cmp437_out0), .out1(cmp437_out1));
cmp cmp438 (.in0(cmp438_in0), .in1(cmp438_in1), .out0(cmp438_out0), .out1(cmp438_out1));
cmp cmp439 (.in0(cmp439_in0), .in1(cmp439_in1), .out0(cmp439_out0), .out1(cmp439_out1));
cmp cmp440 (.in0(cmp440_in0), .in1(cmp440_in1), .out0(cmp440_out0), .out1(cmp440_out1));
cmp cmp441 (.in0(cmp441_in0), .in1(cmp441_in1), .out0(cmp441_out0), .out1(cmp441_out1));
cmp cmp442 (.in0(cmp442_in0), .in1(cmp442_in1), .out0(cmp442_out0), .out1(cmp442_out1));
cmp cmp443 (.in0(cmp443_in0), .in1(cmp443_in1), .out0(cmp443_out0), .out1(cmp443_out1));
cmp cmp444 (.in0(cmp444_in0), .in1(cmp444_in1), .out0(cmp444_out0), .out1(cmp444_out1));
cmp cmp445 (.in0(cmp445_in0), .in1(cmp445_in1), .out0(cmp445_out0), .out1(cmp445_out1));
cmp cmp446 (.in0(cmp446_in0), .in1(cmp446_in1), .out0(cmp446_out0), .out1(cmp446_out1));
cmp cmp447 (.in0(cmp447_in0), .in1(cmp447_in1), .out0(cmp447_out0), .out1(cmp447_out1));
cmp cmp448 (.in0(cmp448_in0), .in1(cmp448_in1), .out0(cmp448_out0), .out1(cmp448_out1));
cmp cmp449 (.in0(cmp449_in0), .in1(cmp449_in1), .out0(cmp449_out0), .out1(cmp449_out1));
cmp cmp450 (.in0(cmp450_in0), .in1(cmp450_in1), .out0(cmp450_out0), .out1(cmp450_out1));
cmp cmp451 (.in0(cmp451_in0), .in1(cmp451_in1), .out0(cmp451_out0), .out1(cmp451_out1));
cmp cmp452 (.in0(cmp452_in0), .in1(cmp452_in1), .out0(cmp452_out0), .out1(cmp452_out1));
cmp cmp453 (.in0(cmp453_in0), .in1(cmp453_in1), .out0(cmp453_out0), .out1(cmp453_out1));
cmp cmp454 (.in0(cmp454_in0), .in1(cmp454_in1), .out0(cmp454_out0), .out1(cmp454_out1));
cmp cmp455 (.in0(cmp455_in0), .in1(cmp455_in1), .out0(cmp455_out0), .out1(cmp455_out1));
cmp cmp456 (.in0(cmp456_in0), .in1(cmp456_in1), .out0(cmp456_out0), .out1(cmp456_out1));
cmp cmp457 (.in0(cmp457_in0), .in1(cmp457_in1), .out0(cmp457_out0), .out1(cmp457_out1));
cmp cmp458 (.in0(cmp458_in0), .in1(cmp458_in1), .out0(cmp458_out0), .out1(cmp458_out1));
cmp cmp459 (.in0(cmp459_in0), .in1(cmp459_in1), .out0(cmp459_out0), .out1(cmp459_out1));
cmp cmp460 (.in0(cmp460_in0), .in1(cmp460_in1), .out0(cmp460_out0), .out1(cmp460_out1));
cmp cmp461 (.in0(cmp461_in0), .in1(cmp461_in1), .out0(cmp461_out0), .out1(cmp461_out1));
cmp cmp462 (.in0(cmp462_in0), .in1(cmp462_in1), .out0(cmp462_out0), .out1(cmp462_out1));
cmp cmp463 (.in0(cmp463_in0), .in1(cmp463_in1), .out0(cmp463_out0), .out1(cmp463_out1));
cmp cmp464 (.in0(cmp464_in0), .in1(cmp464_in1), .out0(cmp464_out0), .out1(cmp464_out1));
cmp cmp465 (.in0(cmp465_in0), .in1(cmp465_in1), .out0(cmp465_out0), .out1(cmp465_out1));
cmp cmp466 (.in0(cmp466_in0), .in1(cmp466_in1), .out0(cmp466_out0), .out1(cmp466_out1));
cmp cmp467 (.in0(cmp467_in0), .in1(cmp467_in1), .out0(cmp467_out0), .out1(cmp467_out1));
cmp cmp468 (.in0(cmp468_in0), .in1(cmp468_in1), .out0(cmp468_out0), .out1(cmp468_out1));
cmp cmp469 (.in0(cmp469_in0), .in1(cmp469_in1), .out0(cmp469_out0), .out1(cmp469_out1));
cmp cmp470 (.in0(cmp470_in0), .in1(cmp470_in1), .out0(cmp470_out0), .out1(cmp470_out1));
cmp cmp471 (.in0(cmp471_in0), .in1(cmp471_in1), .out0(cmp471_out0), .out1(cmp471_out1));
cmp cmp472 (.in0(cmp472_in0), .in1(cmp472_in1), .out0(cmp472_out0), .out1(cmp472_out1));
cmp cmp473 (.in0(cmp473_in0), .in1(cmp473_in1), .out0(cmp473_out0), .out1(cmp473_out1));
cmp cmp474 (.in0(cmp474_in0), .in1(cmp474_in1), .out0(cmp474_out0), .out1(cmp474_out1));
cmp cmp475 (.in0(cmp475_in0), .in1(cmp475_in1), .out0(cmp475_out0), .out1(cmp475_out1));
cmp cmp476 (.in0(cmp476_in0), .in1(cmp476_in1), .out0(cmp476_out0), .out1(cmp476_out1));
cmp cmp477 (.in0(cmp477_in0), .in1(cmp477_in1), .out0(cmp477_out0), .out1(cmp477_out1));
cmp cmp478 (.in0(cmp478_in0), .in1(cmp478_in1), .out0(cmp478_out0), .out1(cmp478_out1));
cmp cmp479 (.in0(cmp479_in0), .in1(cmp479_in1), .out0(cmp479_out0), .out1(cmp479_out1));
cmp cmp480 (.in0(cmp480_in0), .in1(cmp480_in1), .out0(cmp480_out0), .out1(cmp480_out1));
cmp cmp481 (.in0(cmp481_in0), .in1(cmp481_in1), .out0(cmp481_out0), .out1(cmp481_out1));
cmp cmp482 (.in0(cmp482_in0), .in1(cmp482_in1), .out0(cmp482_out0), .out1(cmp482_out1));
cmp cmp483 (.in0(cmp483_in0), .in1(cmp483_in1), .out0(cmp483_out0), .out1(cmp483_out1));
cmp cmp484 (.in0(cmp484_in0), .in1(cmp484_in1), .out0(cmp484_out0), .out1(cmp484_out1));
cmp cmp485 (.in0(cmp485_in0), .in1(cmp485_in1), .out0(cmp485_out0), .out1(cmp485_out1));
cmp cmp486 (.in0(cmp486_in0), .in1(cmp486_in1), .out0(cmp486_out0), .out1(cmp486_out1));
cmp cmp487 (.in0(cmp487_in0), .in1(cmp487_in1), .out0(cmp487_out0), .out1(cmp487_out1));
cmp cmp488 (.in0(cmp488_in0), .in1(cmp488_in1), .out0(cmp488_out0), .out1(cmp488_out1));
cmp cmp489 (.in0(cmp489_in0), .in1(cmp489_in1), .out0(cmp489_out0), .out1(cmp489_out1));
cmp cmp490 (.in0(cmp490_in0), .in1(cmp490_in1), .out0(cmp490_out0), .out1(cmp490_out1));
cmp cmp491 (.in0(cmp491_in0), .in1(cmp491_in1), .out0(cmp491_out0), .out1(cmp491_out1));
cmp cmp492 (.in0(cmp492_in0), .in1(cmp492_in1), .out0(cmp492_out0), .out1(cmp492_out1));
cmp cmp493 (.in0(cmp493_in0), .in1(cmp493_in1), .out0(cmp493_out0), .out1(cmp493_out1));
cmp cmp494 (.in0(cmp494_in0), .in1(cmp494_in1), .out0(cmp494_out0), .out1(cmp494_out1));
cmp cmp495 (.in0(cmp495_in0), .in1(cmp495_in1), .out0(cmp495_out0), .out1(cmp495_out1));
cmp cmp496 (.in0(cmp496_in0), .in1(cmp496_in1), .out0(cmp496_out0), .out1(cmp496_out1));
cmp cmp497 (.in0(cmp497_in0), .in1(cmp497_in1), .out0(cmp497_out0), .out1(cmp497_out1));
cmp cmp498 (.in0(cmp498_in0), .in1(cmp498_in1), .out0(cmp498_out0), .out1(cmp498_out1));
cmp cmp499 (.in0(cmp499_in0), .in1(cmp499_in1), .out0(cmp499_out0), .out1(cmp499_out1));
cmp cmp500 (.in0(cmp500_in0), .in1(cmp500_in1), .out0(cmp500_out0), .out1(cmp500_out1));
cmp cmp501 (.in0(cmp501_in0), .in1(cmp501_in1), .out0(cmp501_out0), .out1(cmp501_out1));
cmp cmp502 (.in0(cmp502_in0), .in1(cmp502_in1), .out0(cmp502_out0), .out1(cmp502_out1));
cmp cmp503 (.in0(cmp503_in0), .in1(cmp503_in1), .out0(cmp503_out0), .out1(cmp503_out1));
cmp cmp504 (.in0(cmp504_in0), .in1(cmp504_in1), .out0(cmp504_out0), .out1(cmp504_out1));
cmp cmp505 (.in0(cmp505_in0), .in1(cmp505_in1), .out0(cmp505_out0), .out1(cmp505_out1));
cmp cmp506 (.in0(cmp506_in0), .in1(cmp506_in1), .out0(cmp506_out0), .out1(cmp506_out1));
cmp cmp507 (.in0(cmp507_in0), .in1(cmp507_in1), .out0(cmp507_out0), .out1(cmp507_out1));
cmp cmp508 (.in0(cmp508_in0), .in1(cmp508_in1), .out0(cmp508_out0), .out1(cmp508_out1));
cmp cmp509 (.in0(cmp509_in0), .in1(cmp509_in1), .out0(cmp509_out0), .out1(cmp509_out1));
cmp cmp510 (.in0(cmp510_in0), .in1(cmp510_in1), .out0(cmp510_out0), .out1(cmp510_out1));
cmp cmp511 (.in0(cmp511_in0), .in1(cmp511_in1), .out0(cmp511_out0), .out1(cmp511_out1));
cmp cmp512 (.in0(cmp512_in0), .in1(cmp512_in1), .out0(cmp512_out0), .out1(cmp512_out1));
cmp cmp513 (.in0(cmp513_in0), .in1(cmp513_in1), .out0(cmp513_out0), .out1(cmp513_out1));
cmp cmp514 (.in0(cmp514_in0), .in1(cmp514_in1), .out0(cmp514_out0), .out1(cmp514_out1));
cmp cmp515 (.in0(cmp515_in0), .in1(cmp515_in1), .out0(cmp515_out0), .out1(cmp515_out1));
cmp cmp516 (.in0(cmp516_in0), .in1(cmp516_in1), .out0(cmp516_out0), .out1(cmp516_out1));
cmp cmp517 (.in0(cmp517_in0), .in1(cmp517_in1), .out0(cmp517_out0), .out1(cmp517_out1));
cmp cmp518 (.in0(cmp518_in0), .in1(cmp518_in1), .out0(cmp518_out0), .out1(cmp518_out1));
cmp cmp519 (.in0(cmp519_in0), .in1(cmp519_in1), .out0(cmp519_out0), .out1(cmp519_out1));
cmp cmp520 (.in0(cmp520_in0), .in1(cmp520_in1), .out0(cmp520_out0), .out1(cmp520_out1));
cmp cmp521 (.in0(cmp521_in0), .in1(cmp521_in1), .out0(cmp521_out0), .out1(cmp521_out1));
cmp cmp522 (.in0(cmp522_in0), .in1(cmp522_in1), .out0(cmp522_out0), .out1(cmp522_out1));
cmp cmp523 (.in0(cmp523_in0), .in1(cmp523_in1), .out0(cmp523_out0), .out1(cmp523_out1));
cmp cmp524 (.in0(cmp524_in0), .in1(cmp524_in1), .out0(cmp524_out0), .out1(cmp524_out1));
cmp cmp525 (.in0(cmp525_in0), .in1(cmp525_in1), .out0(cmp525_out0), .out1(cmp525_out1));
cmp cmp526 (.in0(cmp526_in0), .in1(cmp526_in1), .out0(cmp526_out0), .out1(cmp526_out1));
cmp cmp527 (.in0(cmp527_in0), .in1(cmp527_in1), .out0(cmp527_out0), .out1(cmp527_out1));
cmp cmp528 (.in0(cmp528_in0), .in1(cmp528_in1), .out0(cmp528_out0), .out1(cmp528_out1));
cmp cmp529 (.in0(cmp529_in0), .in1(cmp529_in1), .out0(cmp529_out0), .out1(cmp529_out1));
cmp cmp530 (.in0(cmp530_in0), .in1(cmp530_in1), .out0(cmp530_out0), .out1(cmp530_out1));
cmp cmp531 (.in0(cmp531_in0), .in1(cmp531_in1), .out0(cmp531_out0), .out1(cmp531_out1));
cmp cmp532 (.in0(cmp532_in0), .in1(cmp532_in1), .out0(cmp532_out0), .out1(cmp532_out1));
cmp cmp533 (.in0(cmp533_in0), .in1(cmp533_in1), .out0(cmp533_out0), .out1(cmp533_out1));
cmp cmp534 (.in0(cmp534_in0), .in1(cmp534_in1), .out0(cmp534_out0), .out1(cmp534_out1));
cmp cmp535 (.in0(cmp535_in0), .in1(cmp535_in1), .out0(cmp535_out0), .out1(cmp535_out1));
cmp cmp536 (.in0(cmp536_in0), .in1(cmp536_in1), .out0(cmp536_out0), .out1(cmp536_out1));
cmp cmp537 (.in0(cmp537_in0), .in1(cmp537_in1), .out0(cmp537_out0), .out1(cmp537_out1));
cmp cmp538 (.in0(cmp538_in0), .in1(cmp538_in1), .out0(cmp538_out0), .out1(cmp538_out1));
cmp cmp539 (.in0(cmp539_in0), .in1(cmp539_in1), .out0(cmp539_out0), .out1(cmp539_out1));
cmp cmp540 (.in0(cmp540_in0), .in1(cmp540_in1), .out0(cmp540_out0), .out1(cmp540_out1));
cmp cmp541 (.in0(cmp541_in0), .in1(cmp541_in1), .out0(cmp541_out0), .out1(cmp541_out1));
cmp cmp542 (.in0(cmp542_in0), .in1(cmp542_in1), .out0(cmp542_out0), .out1(cmp542_out1));
cmp cmp543 (.in0(cmp543_in0), .in1(cmp543_in1), .out0(cmp543_out0), .out1(cmp543_out1));
cmp cmp544 (.in0(cmp544_in0), .in1(cmp544_in1), .out0(cmp544_out0), .out1(cmp544_out1));
cmp cmp545 (.in0(cmp545_in0), .in1(cmp545_in1), .out0(cmp545_out0), .out1(cmp545_out1));
cmp cmp546 (.in0(cmp546_in0), .in1(cmp546_in1), .out0(cmp546_out0), .out1(cmp546_out1));
cmp cmp547 (.in0(cmp547_in0), .in1(cmp547_in1), .out0(cmp547_out0), .out1(cmp547_out1));
cmp cmp548 (.in0(cmp548_in0), .in1(cmp548_in1), .out0(cmp548_out0), .out1(cmp548_out1));
cmp cmp549 (.in0(cmp549_in0), .in1(cmp549_in1), .out0(cmp549_out0), .out1(cmp549_out1));
cmp cmp550 (.in0(cmp550_in0), .in1(cmp550_in1), .out0(cmp550_out0), .out1(cmp550_out1));
cmp cmp551 (.in0(cmp551_in0), .in1(cmp551_in1), .out0(cmp551_out0), .out1(cmp551_out1));
cmp cmp552 (.in0(cmp552_in0), .in1(cmp552_in1), .out0(cmp552_out0), .out1(cmp552_out1));
cmp cmp553 (.in0(cmp553_in0), .in1(cmp553_in1), .out0(cmp553_out0), .out1(cmp553_out1));
cmp cmp554 (.in0(cmp554_in0), .in1(cmp554_in1), .out0(cmp554_out0), .out1(cmp554_out1));
cmp cmp555 (.in0(cmp555_in0), .in1(cmp555_in1), .out0(cmp555_out0), .out1(cmp555_out1));
cmp cmp556 (.in0(cmp556_in0), .in1(cmp556_in1), .out0(cmp556_out0), .out1(cmp556_out1));
cmp cmp557 (.in0(cmp557_in0), .in1(cmp557_in1), .out0(cmp557_out0), .out1(cmp557_out1));
cmp cmp558 (.in0(cmp558_in0), .in1(cmp558_in1), .out0(cmp558_out0), .out1(cmp558_out1));
cmp cmp559 (.in0(cmp559_in0), .in1(cmp559_in1), .out0(cmp559_out0), .out1(cmp559_out1));
cmp cmp560 (.in0(cmp560_in0), .in1(cmp560_in1), .out0(cmp560_out0), .out1(cmp560_out1));
cmp cmp561 (.in0(cmp561_in0), .in1(cmp561_in1), .out0(cmp561_out0), .out1(cmp561_out1));
cmp cmp562 (.in0(cmp562_in0), .in1(cmp562_in1), .out0(cmp562_out0), .out1(cmp562_out1));
cmp cmp563 (.in0(cmp563_in0), .in1(cmp563_in1), .out0(cmp563_out0), .out1(cmp563_out1));
cmp cmp564 (.in0(cmp564_in0), .in1(cmp564_in1), .out0(cmp564_out0), .out1(cmp564_out1));
cmp cmp565 (.in0(cmp565_in0), .in1(cmp565_in1), .out0(cmp565_out0), .out1(cmp565_out1));
cmp cmp566 (.in0(cmp566_in0), .in1(cmp566_in1), .out0(cmp566_out0), .out1(cmp566_out1));
cmp cmp567 (.in0(cmp567_in0), .in1(cmp567_in1), .out0(cmp567_out0), .out1(cmp567_out1));
cmp cmp568 (.in0(cmp568_in0), .in1(cmp568_in1), .out0(cmp568_out0), .out1(cmp568_out1));
cmp cmp569 (.in0(cmp569_in0), .in1(cmp569_in1), .out0(cmp569_out0), .out1(cmp569_out1));
cmp cmp570 (.in0(cmp570_in0), .in1(cmp570_in1), .out0(cmp570_out0), .out1(cmp570_out1));
cmp cmp571 (.in0(cmp571_in0), .in1(cmp571_in1), .out0(cmp571_out0), .out1(cmp571_out1));
cmp cmp572 (.in0(cmp572_in0), .in1(cmp572_in1), .out0(cmp572_out0), .out1(cmp572_out1));
cmp cmp573 (.in0(cmp573_in0), .in1(cmp573_in1), .out0(cmp573_out0), .out1(cmp573_out1));
cmp cmp574 (.in0(cmp574_in0), .in1(cmp574_in1), .out0(cmp574_out0), .out1(cmp574_out1));
cmp cmp575 (.in0(cmp575_in0), .in1(cmp575_in1), .out0(cmp575_out0), .out1(cmp575_out1));
cmp cmp576 (.in0(cmp576_in0), .in1(cmp576_in1), .out0(cmp576_out0), .out1(cmp576_out1));
cmp cmp577 (.in0(cmp577_in0), .in1(cmp577_in1), .out0(cmp577_out0), .out1(cmp577_out1));
cmp cmp578 (.in0(cmp578_in0), .in1(cmp578_in1), .out0(cmp578_out0), .out1(cmp578_out1));
cmp cmp579 (.in0(cmp579_in0), .in1(cmp579_in1), .out0(cmp579_out0), .out1(cmp579_out1));
cmp cmp580 (.in0(cmp580_in0), .in1(cmp580_in1), .out0(cmp580_out0), .out1(cmp580_out1));
cmp cmp581 (.in0(cmp581_in0), .in1(cmp581_in1), .out0(cmp581_out0), .out1(cmp581_out1));
cmp cmp582 (.in0(cmp582_in0), .in1(cmp582_in1), .out0(cmp582_out0), .out1(cmp582_out1));
cmp cmp583 (.in0(cmp583_in0), .in1(cmp583_in1), .out0(cmp583_out0), .out1(cmp583_out1));
cmp cmp584 (.in0(cmp584_in0), .in1(cmp584_in1), .out0(cmp584_out0), .out1(cmp584_out1));
cmp cmp585 (.in0(cmp585_in0), .in1(cmp585_in1), .out0(cmp585_out0), .out1(cmp585_out1));
cmp cmp586 (.in0(cmp586_in0), .in1(cmp586_in1), .out0(cmp586_out0), .out1(cmp586_out1));
cmp cmp587 (.in0(cmp587_in0), .in1(cmp587_in1), .out0(cmp587_out0), .out1(cmp587_out1));
cmp cmp588 (.in0(cmp588_in0), .in1(cmp588_in1), .out0(cmp588_out0), .out1(cmp588_out1));
cmp cmp589 (.in0(cmp589_in0), .in1(cmp589_in1), .out0(cmp589_out0), .out1(cmp589_out1));
cmp cmp590 (.in0(cmp590_in0), .in1(cmp590_in1), .out0(cmp590_out0), .out1(cmp590_out1));
cmp cmp591 (.in0(cmp591_in0), .in1(cmp591_in1), .out0(cmp591_out0), .out1(cmp591_out1));
cmp cmp592 (.in0(cmp592_in0), .in1(cmp592_in1), .out0(cmp592_out0), .out1(cmp592_out1));
cmp cmp593 (.in0(cmp593_in0), .in1(cmp593_in1), .out0(cmp593_out0), .out1(cmp593_out1));
cmp cmp594 (.in0(cmp594_in0), .in1(cmp594_in1), .out0(cmp594_out0), .out1(cmp594_out1));
cmp cmp595 (.in0(cmp595_in0), .in1(cmp595_in1), .out0(cmp595_out0), .out1(cmp595_out1));
cmp cmp596 (.in0(cmp596_in0), .in1(cmp596_in1), .out0(cmp596_out0), .out1(cmp596_out1));
cmp cmp597 (.in0(cmp597_in0), .in1(cmp597_in1), .out0(cmp597_out0), .out1(cmp597_out1));
cmp cmp598 (.in0(cmp598_in0), .in1(cmp598_in1), .out0(cmp598_out0), .out1(cmp598_out1));
cmp cmp599 (.in0(cmp599_in0), .in1(cmp599_in1), .out0(cmp599_out0), .out1(cmp599_out1));
cmp cmp600 (.in0(cmp600_in0), .in1(cmp600_in1), .out0(cmp600_out0), .out1(cmp600_out1));
cmp cmp601 (.in0(cmp601_in0), .in1(cmp601_in1), .out0(cmp601_out0), .out1(cmp601_out1));
cmp cmp602 (.in0(cmp602_in0), .in1(cmp602_in1), .out0(cmp602_out0), .out1(cmp602_out1));
cmp cmp603 (.in0(cmp603_in0), .in1(cmp603_in1), .out0(cmp603_out0), .out1(cmp603_out1));
cmp cmp604 (.in0(cmp604_in0), .in1(cmp604_in1), .out0(cmp604_out0), .out1(cmp604_out1));
cmp cmp605 (.in0(cmp605_in0), .in1(cmp605_in1), .out0(cmp605_out0), .out1(cmp605_out1));
cmp cmp606 (.in0(cmp606_in0), .in1(cmp606_in1), .out0(cmp606_out0), .out1(cmp606_out1));
cmp cmp607 (.in0(cmp607_in0), .in1(cmp607_in1), .out0(cmp607_out0), .out1(cmp607_out1));
cmp cmp608 (.in0(cmp608_in0), .in1(cmp608_in1), .out0(cmp608_out0), .out1(cmp608_out1));
cmp cmp609 (.in0(cmp609_in0), .in1(cmp609_in1), .out0(cmp609_out0), .out1(cmp609_out1));
cmp cmp610 (.in0(cmp610_in0), .in1(cmp610_in1), .out0(cmp610_out0), .out1(cmp610_out1));
cmp cmp611 (.in0(cmp611_in0), .in1(cmp611_in1), .out0(cmp611_out0), .out1(cmp611_out1));
cmp cmp612 (.in0(cmp612_in0), .in1(cmp612_in1), .out0(cmp612_out0), .out1(cmp612_out1));
cmp cmp613 (.in0(cmp613_in0), .in1(cmp613_in1), .out0(cmp613_out0), .out1(cmp613_out1));
cmp cmp614 (.in0(cmp614_in0), .in1(cmp614_in1), .out0(cmp614_out0), .out1(cmp614_out1));
cmp cmp615 (.in0(cmp615_in0), .in1(cmp615_in1), .out0(cmp615_out0), .out1(cmp615_out1));
cmp cmp616 (.in0(cmp616_in0), .in1(cmp616_in1), .out0(cmp616_out0), .out1(cmp616_out1));
cmp cmp617 (.in0(cmp617_in0), .in1(cmp617_in1), .out0(cmp617_out0), .out1(cmp617_out1));
cmp cmp618 (.in0(cmp618_in0), .in1(cmp618_in1), .out0(cmp618_out0), .out1(cmp618_out1));
cmp cmp619 (.in0(cmp619_in0), .in1(cmp619_in1), .out0(cmp619_out0), .out1(cmp619_out1));
cmp cmp620 (.in0(cmp620_in0), .in1(cmp620_in1), .out0(cmp620_out0), .out1(cmp620_out1));
cmp cmp621 (.in0(cmp621_in0), .in1(cmp621_in1), .out0(cmp621_out0), .out1(cmp621_out1));
cmp cmp622 (.in0(cmp622_in0), .in1(cmp622_in1), .out0(cmp622_out0), .out1(cmp622_out1));
cmp cmp623 (.in0(cmp623_in0), .in1(cmp623_in1), .out0(cmp623_out0), .out1(cmp623_out1));
cmp cmp624 (.in0(cmp624_in0), .in1(cmp624_in1), .out0(cmp624_out0), .out1(cmp624_out1));
cmp cmp625 (.in0(cmp625_in0), .in1(cmp625_in1), .out0(cmp625_out0), .out1(cmp625_out1));
cmp cmp626 (.in0(cmp626_in0), .in1(cmp626_in1), .out0(cmp626_out0), .out1(cmp626_out1));
cmp cmp627 (.in0(cmp627_in0), .in1(cmp627_in1), .out0(cmp627_out0), .out1(cmp627_out1));
cmp cmp628 (.in0(cmp628_in0), .in1(cmp628_in1), .out0(cmp628_out0), .out1(cmp628_out1));
cmp cmp629 (.in0(cmp629_in0), .in1(cmp629_in1), .out0(cmp629_out0), .out1(cmp629_out1));
cmp cmp630 (.in0(cmp630_in0), .in1(cmp630_in1), .out0(cmp630_out0), .out1(cmp630_out1));
cmp cmp631 (.in0(cmp631_in0), .in1(cmp631_in1), .out0(cmp631_out0), .out1(cmp631_out1));
cmp cmp632 (.in0(cmp632_in0), .in1(cmp632_in1), .out0(cmp632_out0), .out1(cmp632_out1));
cmp cmp633 (.in0(cmp633_in0), .in1(cmp633_in1), .out0(cmp633_out0), .out1(cmp633_out1));
cmp cmp634 (.in0(cmp634_in0), .in1(cmp634_in1), .out0(cmp634_out0), .out1(cmp634_out1));
cmp cmp635 (.in0(cmp635_in0), .in1(cmp635_in1), .out0(cmp635_out0), .out1(cmp635_out1));
cmp cmp636 (.in0(cmp636_in0), .in1(cmp636_in1), .out0(cmp636_out0), .out1(cmp636_out1));
cmp cmp637 (.in0(cmp637_in0), .in1(cmp637_in1), .out0(cmp637_out0), .out1(cmp637_out1));
cmp cmp638 (.in0(cmp638_in0), .in1(cmp638_in1), .out0(cmp638_out0), .out1(cmp638_out1));
cmp cmp639 (.in0(cmp639_in0), .in1(cmp639_in1), .out0(cmp639_out0), .out1(cmp639_out1));
cmp cmp640 (.in0(cmp640_in0), .in1(cmp640_in1), .out0(cmp640_out0), .out1(cmp640_out1));
cmp cmp641 (.in0(cmp641_in0), .in1(cmp641_in1), .out0(cmp641_out0), .out1(cmp641_out1));
cmp cmp642 (.in0(cmp642_in0), .in1(cmp642_in1), .out0(cmp642_out0), .out1(cmp642_out1));
cmp cmp643 (.in0(cmp643_in0), .in1(cmp643_in1), .out0(cmp643_out0), .out1(cmp643_out1));
cmp cmp644 (.in0(cmp644_in0), .in1(cmp644_in1), .out0(cmp644_out0), .out1(cmp644_out1));
cmp cmp645 (.in0(cmp645_in0), .in1(cmp645_in1), .out0(cmp645_out0), .out1(cmp645_out1));
cmp cmp646 (.in0(cmp646_in0), .in1(cmp646_in1), .out0(cmp646_out0), .out1(cmp646_out1));
cmp cmp647 (.in0(cmp647_in0), .in1(cmp647_in1), .out0(cmp647_out0), .out1(cmp647_out1));
cmp cmp648 (.in0(cmp648_in0), .in1(cmp648_in1), .out0(cmp648_out0), .out1(cmp648_out1));
cmp cmp649 (.in0(cmp649_in0), .in1(cmp649_in1), .out0(cmp649_out0), .out1(cmp649_out1));
cmp cmp650 (.in0(cmp650_in0), .in1(cmp650_in1), .out0(cmp650_out0), .out1(cmp650_out1));
cmp cmp651 (.in0(cmp651_in0), .in1(cmp651_in1), .out0(cmp651_out0), .out1(cmp651_out1));
cmp cmp652 (.in0(cmp652_in0), .in1(cmp652_in1), .out0(cmp652_out0), .out1(cmp652_out1));
cmp cmp653 (.in0(cmp653_in0), .in1(cmp653_in1), .out0(cmp653_out0), .out1(cmp653_out1));
cmp cmp654 (.in0(cmp654_in0), .in1(cmp654_in1), .out0(cmp654_out0), .out1(cmp654_out1));
cmp cmp655 (.in0(cmp655_in0), .in1(cmp655_in1), .out0(cmp655_out0), .out1(cmp655_out1));
cmp cmp656 (.in0(cmp656_in0), .in1(cmp656_in1), .out0(cmp656_out0), .out1(cmp656_out1));
cmp cmp657 (.in0(cmp657_in0), .in1(cmp657_in1), .out0(cmp657_out0), .out1(cmp657_out1));
cmp cmp658 (.in0(cmp658_in0), .in1(cmp658_in1), .out0(cmp658_out0), .out1(cmp658_out1));
cmp cmp659 (.in0(cmp659_in0), .in1(cmp659_in1), .out0(cmp659_out0), .out1(cmp659_out1));
cmp cmp660 (.in0(cmp660_in0), .in1(cmp660_in1), .out0(cmp660_out0), .out1(cmp660_out1));
assign median = cmp660_out1;
endmodule

//--------------comparator----------------
module cmp(
     input  [7:0] in0,
     input  [7:0] in1,
     output wire [7:0] out0,
     output wire [7:0] out1
);
     assign out0 = (in0<in1) ? in0:in1;
     assign out1 = (in0<in1) ? in1:in0;
endmodule
